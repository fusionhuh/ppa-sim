`ifndef CARRY_OPERATOR
`include "carry_operator.v"
`endif
`ifndef NEG_CARRY_OPERATOR
`include "neg_operator.v"
`endif
`ifndef POS_CARRY_OPERATOR
`include "pos_operator.v"
`endif
// number of levels: 11
// number of nodes: 253
module hybridadder128_4(x1, x2, s);
	input[127:0]x1;
	input[127:0]x2;
	output[127:0]s;
	wire[127:0]p_in = x1 ^ x2;
	wire[127:0]g_in = x1 & x2;
	wire node_level1_pos1_outg;
	wire node_level1_pos1_outp;
	neg_operator node_level1_pos1(.p1(p_in[1]), .g1(g_in[1]), .p0(p_in[0]), .g0(g_in[0]), .gp(node_level1_pos1_outg), .pp(node_level1_pos1_outp));
	wire node_level1_pos3_outg;
	wire node_level1_pos3_outp;
	neg_operator node_level1_pos3(.p1(p_in[3]), .g1(g_in[3]), .p0(p_in[2]), .g0(g_in[2]), .gp(node_level1_pos3_outg), .pp(node_level1_pos3_outp));
	wire node_level1_pos5_outg;
	wire node_level1_pos5_outp;
	neg_operator node_level1_pos5(.p1(p_in[5]), .g1(g_in[5]), .p0(p_in[4]), .g0(g_in[4]), .gp(node_level1_pos5_outg), .pp(node_level1_pos5_outp));
	wire node_level1_pos7_outg;
	wire node_level1_pos7_outp;
	neg_operator node_level1_pos7(.p1(p_in[7]), .g1(g_in[7]), .p0(p_in[6]), .g0(g_in[6]), .gp(node_level1_pos7_outg), .pp(node_level1_pos7_outp));
	wire node_level1_pos9_outg;
	wire node_level1_pos9_outp;
	neg_operator node_level1_pos9(.p1(p_in[9]), .g1(g_in[9]), .p0(p_in[8]), .g0(g_in[8]), .gp(node_level1_pos9_outg), .pp(node_level1_pos9_outp));
	wire node_level1_pos11_outg;
	wire node_level1_pos11_outp;
	neg_operator node_level1_pos11(.p1(p_in[11]), .g1(g_in[11]), .p0(p_in[10]), .g0(g_in[10]), .gp(node_level1_pos11_outg), .pp(node_level1_pos11_outp));
	wire node_level1_pos13_outg;
	wire node_level1_pos13_outp;
	neg_operator node_level1_pos13(.p1(p_in[13]), .g1(g_in[13]), .p0(p_in[12]), .g0(g_in[12]), .gp(node_level1_pos13_outg), .pp(node_level1_pos13_outp));
	wire node_level1_pos15_outg;
	wire node_level1_pos15_outp;
	neg_operator node_level1_pos15(.p1(p_in[15]), .g1(g_in[15]), .p0(p_in[14]), .g0(g_in[14]), .gp(node_level1_pos15_outg), .pp(node_level1_pos15_outp));
	wire node_level1_pos17_outg;
	wire node_level1_pos17_outp;
	neg_operator node_level1_pos17(.p1(p_in[17]), .g1(g_in[17]), .p0(p_in[16]), .g0(g_in[16]), .gp(node_level1_pos17_outg), .pp(node_level1_pos17_outp));
	wire node_level1_pos19_outg;
	wire node_level1_pos19_outp;
	neg_operator node_level1_pos19(.p1(p_in[19]), .g1(g_in[19]), .p0(p_in[18]), .g0(g_in[18]), .gp(node_level1_pos19_outg), .pp(node_level1_pos19_outp));
	wire node_level1_pos21_outg;
	wire node_level1_pos21_outp;
	neg_operator node_level1_pos21(.p1(p_in[21]), .g1(g_in[21]), .p0(p_in[20]), .g0(g_in[20]), .gp(node_level1_pos21_outg), .pp(node_level1_pos21_outp));
	wire node_level1_pos23_outg;
	wire node_level1_pos23_outp;
	neg_operator node_level1_pos23(.p1(p_in[23]), .g1(g_in[23]), .p0(p_in[22]), .g0(g_in[22]), .gp(node_level1_pos23_outg), .pp(node_level1_pos23_outp));
	wire node_level1_pos25_outg;
	wire node_level1_pos25_outp;
	neg_operator node_level1_pos25(.p1(p_in[25]), .g1(g_in[25]), .p0(p_in[24]), .g0(g_in[24]), .gp(node_level1_pos25_outg), .pp(node_level1_pos25_outp));
	wire node_level1_pos27_outg;
	wire node_level1_pos27_outp;
	neg_operator node_level1_pos27(.p1(p_in[27]), .g1(g_in[27]), .p0(p_in[26]), .g0(g_in[26]), .gp(node_level1_pos27_outg), .pp(node_level1_pos27_outp));
	wire node_level1_pos29_outg;
	wire node_level1_pos29_outp;
	neg_operator node_level1_pos29(.p1(p_in[29]), .g1(g_in[29]), .p0(p_in[28]), .g0(g_in[28]), .gp(node_level1_pos29_outg), .pp(node_level1_pos29_outp));
	wire node_level1_pos31_outg;
	wire node_level1_pos31_outp;
	neg_operator node_level1_pos31(.p1(p_in[31]), .g1(g_in[31]), .p0(p_in[30]), .g0(g_in[30]), .gp(node_level1_pos31_outg), .pp(node_level1_pos31_outp));
	wire node_level1_pos33_outg;
	wire node_level1_pos33_outp;
	neg_operator node_level1_pos33(.p1(p_in[33]), .g1(g_in[33]), .p0(p_in[32]), .g0(g_in[32]), .gp(node_level1_pos33_outg), .pp(node_level1_pos33_outp));
	wire node_level1_pos35_outg;
	wire node_level1_pos35_outp;
	neg_operator node_level1_pos35(.p1(p_in[35]), .g1(g_in[35]), .p0(p_in[34]), .g0(g_in[34]), .gp(node_level1_pos35_outg), .pp(node_level1_pos35_outp));
	wire node_level1_pos37_outg;
	wire node_level1_pos37_outp;
	neg_operator node_level1_pos37(.p1(p_in[37]), .g1(g_in[37]), .p0(p_in[36]), .g0(g_in[36]), .gp(node_level1_pos37_outg), .pp(node_level1_pos37_outp));
	wire node_level1_pos39_outg;
	wire node_level1_pos39_outp;
	neg_operator node_level1_pos39(.p1(p_in[39]), .g1(g_in[39]), .p0(p_in[38]), .g0(g_in[38]), .gp(node_level1_pos39_outg), .pp(node_level1_pos39_outp));
	wire node_level1_pos41_outg;
	wire node_level1_pos41_outp;
	neg_operator node_level1_pos41(.p1(p_in[41]), .g1(g_in[41]), .p0(p_in[40]), .g0(g_in[40]), .gp(node_level1_pos41_outg), .pp(node_level1_pos41_outp));
	wire node_level1_pos43_outg;
	wire node_level1_pos43_outp;
	neg_operator node_level1_pos43(.p1(p_in[43]), .g1(g_in[43]), .p0(p_in[42]), .g0(g_in[42]), .gp(node_level1_pos43_outg), .pp(node_level1_pos43_outp));
	wire node_level1_pos45_outg;
	wire node_level1_pos45_outp;
	neg_operator node_level1_pos45(.p1(p_in[45]), .g1(g_in[45]), .p0(p_in[44]), .g0(g_in[44]), .gp(node_level1_pos45_outg), .pp(node_level1_pos45_outp));
	wire node_level1_pos47_outg;
	wire node_level1_pos47_outp;
	neg_operator node_level1_pos47(.p1(p_in[47]), .g1(g_in[47]), .p0(p_in[46]), .g0(g_in[46]), .gp(node_level1_pos47_outg), .pp(node_level1_pos47_outp));
	wire node_level1_pos49_outg;
	wire node_level1_pos49_outp;
	neg_operator node_level1_pos49(.p1(p_in[49]), .g1(g_in[49]), .p0(p_in[48]), .g0(g_in[48]), .gp(node_level1_pos49_outg), .pp(node_level1_pos49_outp));
	wire node_level1_pos51_outg;
	wire node_level1_pos51_outp;
	neg_operator node_level1_pos51(.p1(p_in[51]), .g1(g_in[51]), .p0(p_in[50]), .g0(g_in[50]), .gp(node_level1_pos51_outg), .pp(node_level1_pos51_outp));
	wire node_level1_pos53_outg;
	wire node_level1_pos53_outp;
	neg_operator node_level1_pos53(.p1(p_in[53]), .g1(g_in[53]), .p0(p_in[52]), .g0(g_in[52]), .gp(node_level1_pos53_outg), .pp(node_level1_pos53_outp));
	wire node_level1_pos55_outg;
	wire node_level1_pos55_outp;
	neg_operator node_level1_pos55(.p1(p_in[55]), .g1(g_in[55]), .p0(p_in[54]), .g0(g_in[54]), .gp(node_level1_pos55_outg), .pp(node_level1_pos55_outp));
	wire node_level1_pos57_outg;
	wire node_level1_pos57_outp;
	neg_operator node_level1_pos57(.p1(p_in[57]), .g1(g_in[57]), .p0(p_in[56]), .g0(g_in[56]), .gp(node_level1_pos57_outg), .pp(node_level1_pos57_outp));
	wire node_level1_pos59_outg;
	wire node_level1_pos59_outp;
	neg_operator node_level1_pos59(.p1(p_in[59]), .g1(g_in[59]), .p0(p_in[58]), .g0(g_in[58]), .gp(node_level1_pos59_outg), .pp(node_level1_pos59_outp));
	wire node_level1_pos61_outg;
	wire node_level1_pos61_outp;
	neg_operator node_level1_pos61(.p1(p_in[61]), .g1(g_in[61]), .p0(p_in[60]), .g0(g_in[60]), .gp(node_level1_pos61_outg), .pp(node_level1_pos61_outp));
	wire node_level1_pos63_outg;
	wire node_level1_pos63_outp;
	neg_operator node_level1_pos63(.p1(p_in[63]), .g1(g_in[63]), .p0(p_in[62]), .g0(g_in[62]), .gp(node_level1_pos63_outg), .pp(node_level1_pos63_outp));
	wire node_level1_pos65_outg;
	wire node_level1_pos65_outp;
	neg_operator node_level1_pos65(.p1(p_in[65]), .g1(g_in[65]), .p0(p_in[64]), .g0(g_in[64]), .gp(node_level1_pos65_outg), .pp(node_level1_pos65_outp));
	wire node_level1_pos67_outg;
	wire node_level1_pos67_outp;
	neg_operator node_level1_pos67(.p1(p_in[67]), .g1(g_in[67]), .p0(p_in[66]), .g0(g_in[66]), .gp(node_level1_pos67_outg), .pp(node_level1_pos67_outp));
	wire node_level1_pos69_outg;
	wire node_level1_pos69_outp;
	neg_operator node_level1_pos69(.p1(p_in[69]), .g1(g_in[69]), .p0(p_in[68]), .g0(g_in[68]), .gp(node_level1_pos69_outg), .pp(node_level1_pos69_outp));
	wire node_level1_pos71_outg;
	wire node_level1_pos71_outp;
	neg_operator node_level1_pos71(.p1(p_in[71]), .g1(g_in[71]), .p0(p_in[70]), .g0(g_in[70]), .gp(node_level1_pos71_outg), .pp(node_level1_pos71_outp));
	wire node_level1_pos73_outg;
	wire node_level1_pos73_outp;
	neg_operator node_level1_pos73(.p1(p_in[73]), .g1(g_in[73]), .p0(p_in[72]), .g0(g_in[72]), .gp(node_level1_pos73_outg), .pp(node_level1_pos73_outp));
	wire node_level1_pos75_outg;
	wire node_level1_pos75_outp;
	neg_operator node_level1_pos75(.p1(p_in[75]), .g1(g_in[75]), .p0(p_in[74]), .g0(g_in[74]), .gp(node_level1_pos75_outg), .pp(node_level1_pos75_outp));
	wire node_level1_pos77_outg;
	wire node_level1_pos77_outp;
	neg_operator node_level1_pos77(.p1(p_in[77]), .g1(g_in[77]), .p0(p_in[76]), .g0(g_in[76]), .gp(node_level1_pos77_outg), .pp(node_level1_pos77_outp));
	wire node_level1_pos79_outg;
	wire node_level1_pos79_outp;
	neg_operator node_level1_pos79(.p1(p_in[79]), .g1(g_in[79]), .p0(p_in[78]), .g0(g_in[78]), .gp(node_level1_pos79_outg), .pp(node_level1_pos79_outp));
	wire node_level1_pos81_outg;
	wire node_level1_pos81_outp;
	neg_operator node_level1_pos81(.p1(p_in[81]), .g1(g_in[81]), .p0(p_in[80]), .g0(g_in[80]), .gp(node_level1_pos81_outg), .pp(node_level1_pos81_outp));
	wire node_level1_pos83_outg;
	wire node_level1_pos83_outp;
	neg_operator node_level1_pos83(.p1(p_in[83]), .g1(g_in[83]), .p0(p_in[82]), .g0(g_in[82]), .gp(node_level1_pos83_outg), .pp(node_level1_pos83_outp));
	wire node_level1_pos85_outg;
	wire node_level1_pos85_outp;
	neg_operator node_level1_pos85(.p1(p_in[85]), .g1(g_in[85]), .p0(p_in[84]), .g0(g_in[84]), .gp(node_level1_pos85_outg), .pp(node_level1_pos85_outp));
	wire node_level1_pos87_outg;
	wire node_level1_pos87_outp;
	neg_operator node_level1_pos87(.p1(p_in[87]), .g1(g_in[87]), .p0(p_in[86]), .g0(g_in[86]), .gp(node_level1_pos87_outg), .pp(node_level1_pos87_outp));
	wire node_level1_pos89_outg;
	wire node_level1_pos89_outp;
	neg_operator node_level1_pos89(.p1(p_in[89]), .g1(g_in[89]), .p0(p_in[88]), .g0(g_in[88]), .gp(node_level1_pos89_outg), .pp(node_level1_pos89_outp));
	wire node_level1_pos91_outg;
	wire node_level1_pos91_outp;
	neg_operator node_level1_pos91(.p1(p_in[91]), .g1(g_in[91]), .p0(p_in[90]), .g0(g_in[90]), .gp(node_level1_pos91_outg), .pp(node_level1_pos91_outp));
	wire node_level1_pos93_outg;
	wire node_level1_pos93_outp;
	neg_operator node_level1_pos93(.p1(p_in[93]), .g1(g_in[93]), .p0(p_in[92]), .g0(g_in[92]), .gp(node_level1_pos93_outg), .pp(node_level1_pos93_outp));
	wire node_level1_pos95_outg;
	wire node_level1_pos95_outp;
	neg_operator node_level1_pos95(.p1(p_in[95]), .g1(g_in[95]), .p0(p_in[94]), .g0(g_in[94]), .gp(node_level1_pos95_outg), .pp(node_level1_pos95_outp));
	wire node_level1_pos97_outg;
	wire node_level1_pos97_outp;
	neg_operator node_level1_pos97(.p1(p_in[97]), .g1(g_in[97]), .p0(p_in[96]), .g0(g_in[96]), .gp(node_level1_pos97_outg), .pp(node_level1_pos97_outp));
	wire node_level1_pos99_outg;
	wire node_level1_pos99_outp;
	neg_operator node_level1_pos99(.p1(p_in[99]), .g1(g_in[99]), .p0(p_in[98]), .g0(g_in[98]), .gp(node_level1_pos99_outg), .pp(node_level1_pos99_outp));
	wire node_level1_pos101_outg;
	wire node_level1_pos101_outp;
	neg_operator node_level1_pos101(.p1(p_in[101]), .g1(g_in[101]), .p0(p_in[100]), .g0(g_in[100]), .gp(node_level1_pos101_outg), .pp(node_level1_pos101_outp));
	wire node_level1_pos103_outg;
	wire node_level1_pos103_outp;
	neg_operator node_level1_pos103(.p1(p_in[103]), .g1(g_in[103]), .p0(p_in[102]), .g0(g_in[102]), .gp(node_level1_pos103_outg), .pp(node_level1_pos103_outp));
	wire node_level1_pos105_outg;
	wire node_level1_pos105_outp;
	neg_operator node_level1_pos105(.p1(p_in[105]), .g1(g_in[105]), .p0(p_in[104]), .g0(g_in[104]), .gp(node_level1_pos105_outg), .pp(node_level1_pos105_outp));
	wire node_level1_pos107_outg;
	wire node_level1_pos107_outp;
	neg_operator node_level1_pos107(.p1(p_in[107]), .g1(g_in[107]), .p0(p_in[106]), .g0(g_in[106]), .gp(node_level1_pos107_outg), .pp(node_level1_pos107_outp));
	wire node_level1_pos109_outg;
	wire node_level1_pos109_outp;
	neg_operator node_level1_pos109(.p1(p_in[109]), .g1(g_in[109]), .p0(p_in[108]), .g0(g_in[108]), .gp(node_level1_pos109_outg), .pp(node_level1_pos109_outp));
	wire node_level1_pos111_outg;
	wire node_level1_pos111_outp;
	neg_operator node_level1_pos111(.p1(p_in[111]), .g1(g_in[111]), .p0(p_in[110]), .g0(g_in[110]), .gp(node_level1_pos111_outg), .pp(node_level1_pos111_outp));
	wire node_level1_pos113_outg;
	wire node_level1_pos113_outp;
	neg_operator node_level1_pos113(.p1(p_in[113]), .g1(g_in[113]), .p0(p_in[112]), .g0(g_in[112]), .gp(node_level1_pos113_outg), .pp(node_level1_pos113_outp));
	wire node_level1_pos115_outg;
	wire node_level1_pos115_outp;
	neg_operator node_level1_pos115(.p1(p_in[115]), .g1(g_in[115]), .p0(p_in[114]), .g0(g_in[114]), .gp(node_level1_pos115_outg), .pp(node_level1_pos115_outp));
	wire node_level1_pos117_outg;
	wire node_level1_pos117_outp;
	neg_operator node_level1_pos117(.p1(p_in[117]), .g1(g_in[117]), .p0(p_in[116]), .g0(g_in[116]), .gp(node_level1_pos117_outg), .pp(node_level1_pos117_outp));
	wire node_level1_pos119_outg;
	wire node_level1_pos119_outp;
	neg_operator node_level1_pos119(.p1(p_in[119]), .g1(g_in[119]), .p0(p_in[118]), .g0(g_in[118]), .gp(node_level1_pos119_outg), .pp(node_level1_pos119_outp));
	wire node_level1_pos121_outg;
	wire node_level1_pos121_outp;
	neg_operator node_level1_pos121(.p1(p_in[121]), .g1(g_in[121]), .p0(p_in[120]), .g0(g_in[120]), .gp(node_level1_pos121_outg), .pp(node_level1_pos121_outp));
	wire node_level1_pos123_outg;
	wire node_level1_pos123_outp;
	neg_operator node_level1_pos123(.p1(p_in[123]), .g1(g_in[123]), .p0(p_in[122]), .g0(g_in[122]), .gp(node_level1_pos123_outg), .pp(node_level1_pos123_outp));
	wire node_level1_pos125_outg;
	wire node_level1_pos125_outp;
	neg_operator node_level1_pos125(.p1(p_in[125]), .g1(g_in[125]), .p0(p_in[124]), .g0(g_in[124]), .gp(node_level1_pos125_outg), .pp(node_level1_pos125_outp));
	wire node_level1_pos127_outg;
	wire node_level1_pos127_outp;
	neg_operator node_level1_pos127(.p1(p_in[127]), .g1(g_in[127]), .p0(p_in[126]), .g0(g_in[126]), .gp(node_level1_pos127_outg), .pp(node_level1_pos127_outp));
	wire node_level2_pos3_outg;
	wire node_level2_pos3_outp;
	pos_operator node_level2_pos3(.p1(node_level1_pos3_outp), .g1(node_level1_pos3_outg), .p0(node_level1_pos1_outp), .g0(node_level1_pos1_outg), .gp(node_level2_pos3_outg), .pp(node_level2_pos3_outp));
	wire node_level2_pos7_outg;
	wire node_level2_pos7_outp;
	pos_operator node_level2_pos7(.p1(node_level1_pos7_outp), .g1(node_level1_pos7_outg), .p0(node_level1_pos5_outp), .g0(node_level1_pos5_outg), .gp(node_level2_pos7_outg), .pp(node_level2_pos7_outp));
	wire node_level2_pos11_outg;
	wire node_level2_pos11_outp;
	pos_operator node_level2_pos11(.p1(node_level1_pos11_outp), .g1(node_level1_pos11_outg), .p0(node_level1_pos9_outp), .g0(node_level1_pos9_outg), .gp(node_level2_pos11_outg), .pp(node_level2_pos11_outp));
	wire node_level2_pos15_outg;
	wire node_level2_pos15_outp;
	pos_operator node_level2_pos15(.p1(node_level1_pos15_outp), .g1(node_level1_pos15_outg), .p0(node_level1_pos13_outp), .g0(node_level1_pos13_outg), .gp(node_level2_pos15_outg), .pp(node_level2_pos15_outp));
	wire node_level2_pos19_outg;
	wire node_level2_pos19_outp;
	pos_operator node_level2_pos19(.p1(node_level1_pos19_outp), .g1(node_level1_pos19_outg), .p0(node_level1_pos17_outp), .g0(node_level1_pos17_outg), .gp(node_level2_pos19_outg), .pp(node_level2_pos19_outp));
	wire node_level2_pos23_outg;
	wire node_level2_pos23_outp;
	pos_operator node_level2_pos23(.p1(node_level1_pos23_outp), .g1(node_level1_pos23_outg), .p0(node_level1_pos21_outp), .g0(node_level1_pos21_outg), .gp(node_level2_pos23_outg), .pp(node_level2_pos23_outp));
	wire node_level2_pos27_outg;
	wire node_level2_pos27_outp;
	pos_operator node_level2_pos27(.p1(node_level1_pos27_outp), .g1(node_level1_pos27_outg), .p0(node_level1_pos25_outp), .g0(node_level1_pos25_outg), .gp(node_level2_pos27_outg), .pp(node_level2_pos27_outp));
	wire node_level2_pos31_outg;
	wire node_level2_pos31_outp;
	pos_operator node_level2_pos31(.p1(node_level1_pos31_outp), .g1(node_level1_pos31_outg), .p0(node_level1_pos29_outp), .g0(node_level1_pos29_outg), .gp(node_level2_pos31_outg), .pp(node_level2_pos31_outp));
	wire node_level2_pos35_outg;
	wire node_level2_pos35_outp;
	pos_operator node_level2_pos35(.p1(node_level1_pos35_outp), .g1(node_level1_pos35_outg), .p0(node_level1_pos33_outp), .g0(node_level1_pos33_outg), .gp(node_level2_pos35_outg), .pp(node_level2_pos35_outp));
	wire node_level2_pos39_outg;
	wire node_level2_pos39_outp;
	pos_operator node_level2_pos39(.p1(node_level1_pos39_outp), .g1(node_level1_pos39_outg), .p0(node_level1_pos37_outp), .g0(node_level1_pos37_outg), .gp(node_level2_pos39_outg), .pp(node_level2_pos39_outp));
	wire node_level2_pos43_outg;
	wire node_level2_pos43_outp;
	pos_operator node_level2_pos43(.p1(node_level1_pos43_outp), .g1(node_level1_pos43_outg), .p0(node_level1_pos41_outp), .g0(node_level1_pos41_outg), .gp(node_level2_pos43_outg), .pp(node_level2_pos43_outp));
	wire node_level2_pos47_outg;
	wire node_level2_pos47_outp;
	pos_operator node_level2_pos47(.p1(node_level1_pos47_outp), .g1(node_level1_pos47_outg), .p0(node_level1_pos45_outp), .g0(node_level1_pos45_outg), .gp(node_level2_pos47_outg), .pp(node_level2_pos47_outp));
	wire node_level2_pos51_outg;
	wire node_level2_pos51_outp;
	pos_operator node_level2_pos51(.p1(node_level1_pos51_outp), .g1(node_level1_pos51_outg), .p0(node_level1_pos49_outp), .g0(node_level1_pos49_outg), .gp(node_level2_pos51_outg), .pp(node_level2_pos51_outp));
	wire node_level2_pos55_outg;
	wire node_level2_pos55_outp;
	pos_operator node_level2_pos55(.p1(node_level1_pos55_outp), .g1(node_level1_pos55_outg), .p0(node_level1_pos53_outp), .g0(node_level1_pos53_outg), .gp(node_level2_pos55_outg), .pp(node_level2_pos55_outp));
	wire node_level2_pos59_outg;
	wire node_level2_pos59_outp;
	pos_operator node_level2_pos59(.p1(node_level1_pos59_outp), .g1(node_level1_pos59_outg), .p0(node_level1_pos57_outp), .g0(node_level1_pos57_outg), .gp(node_level2_pos59_outg), .pp(node_level2_pos59_outp));
	wire node_level2_pos63_outg;
	wire node_level2_pos63_outp;
	pos_operator node_level2_pos63(.p1(node_level1_pos63_outp), .g1(node_level1_pos63_outg), .p0(node_level1_pos61_outp), .g0(node_level1_pos61_outg), .gp(node_level2_pos63_outg), .pp(node_level2_pos63_outp));
	wire node_level2_pos67_outg;
	wire node_level2_pos67_outp;
	pos_operator node_level2_pos67(.p1(node_level1_pos67_outp), .g1(node_level1_pos67_outg), .p0(node_level1_pos65_outp), .g0(node_level1_pos65_outg), .gp(node_level2_pos67_outg), .pp(node_level2_pos67_outp));
	wire node_level2_pos71_outg;
	wire node_level2_pos71_outp;
	pos_operator node_level2_pos71(.p1(node_level1_pos71_outp), .g1(node_level1_pos71_outg), .p0(node_level1_pos69_outp), .g0(node_level1_pos69_outg), .gp(node_level2_pos71_outg), .pp(node_level2_pos71_outp));
	wire node_level2_pos75_outg;
	wire node_level2_pos75_outp;
	pos_operator node_level2_pos75(.p1(node_level1_pos75_outp), .g1(node_level1_pos75_outg), .p0(node_level1_pos73_outp), .g0(node_level1_pos73_outg), .gp(node_level2_pos75_outg), .pp(node_level2_pos75_outp));
	wire node_level2_pos79_outg;
	wire node_level2_pos79_outp;
	pos_operator node_level2_pos79(.p1(node_level1_pos79_outp), .g1(node_level1_pos79_outg), .p0(node_level1_pos77_outp), .g0(node_level1_pos77_outg), .gp(node_level2_pos79_outg), .pp(node_level2_pos79_outp));
	wire node_level2_pos83_outg;
	wire node_level2_pos83_outp;
	pos_operator node_level2_pos83(.p1(node_level1_pos83_outp), .g1(node_level1_pos83_outg), .p0(node_level1_pos81_outp), .g0(node_level1_pos81_outg), .gp(node_level2_pos83_outg), .pp(node_level2_pos83_outp));
	wire node_level2_pos87_outg;
	wire node_level2_pos87_outp;
	pos_operator node_level2_pos87(.p1(node_level1_pos87_outp), .g1(node_level1_pos87_outg), .p0(node_level1_pos85_outp), .g0(node_level1_pos85_outg), .gp(node_level2_pos87_outg), .pp(node_level2_pos87_outp));
	wire node_level2_pos91_outg;
	wire node_level2_pos91_outp;
	pos_operator node_level2_pos91(.p1(node_level1_pos91_outp), .g1(node_level1_pos91_outg), .p0(node_level1_pos89_outp), .g0(node_level1_pos89_outg), .gp(node_level2_pos91_outg), .pp(node_level2_pos91_outp));
	wire node_level2_pos95_outg;
	wire node_level2_pos95_outp;
	pos_operator node_level2_pos95(.p1(node_level1_pos95_outp), .g1(node_level1_pos95_outg), .p0(node_level1_pos93_outp), .g0(node_level1_pos93_outg), .gp(node_level2_pos95_outg), .pp(node_level2_pos95_outp));
	wire node_level2_pos99_outg;
	wire node_level2_pos99_outp;
	pos_operator node_level2_pos99(.p1(node_level1_pos99_outp), .g1(node_level1_pos99_outg), .p0(node_level1_pos97_outp), .g0(node_level1_pos97_outg), .gp(node_level2_pos99_outg), .pp(node_level2_pos99_outp));
	wire node_level2_pos103_outg;
	wire node_level2_pos103_outp;
	pos_operator node_level2_pos103(.p1(node_level1_pos103_outp), .g1(node_level1_pos103_outg), .p0(node_level1_pos101_outp), .g0(node_level1_pos101_outg), .gp(node_level2_pos103_outg), .pp(node_level2_pos103_outp));
	wire node_level2_pos107_outg;
	wire node_level2_pos107_outp;
	pos_operator node_level2_pos107(.p1(node_level1_pos107_outp), .g1(node_level1_pos107_outg), .p0(node_level1_pos105_outp), .g0(node_level1_pos105_outg), .gp(node_level2_pos107_outg), .pp(node_level2_pos107_outp));
	wire node_level2_pos111_outg;
	wire node_level2_pos111_outp;
	pos_operator node_level2_pos111(.p1(node_level1_pos111_outp), .g1(node_level1_pos111_outg), .p0(node_level1_pos109_outp), .g0(node_level1_pos109_outg), .gp(node_level2_pos111_outg), .pp(node_level2_pos111_outp));
	wire node_level2_pos115_outg;
	wire node_level2_pos115_outp;
	pos_operator node_level2_pos115(.p1(node_level1_pos115_outp), .g1(node_level1_pos115_outg), .p0(node_level1_pos113_outp), .g0(node_level1_pos113_outg), .gp(node_level2_pos115_outg), .pp(node_level2_pos115_outp));
	wire node_level2_pos119_outg;
	wire node_level2_pos119_outp;
	pos_operator node_level2_pos119(.p1(node_level1_pos119_outp), .g1(node_level1_pos119_outg), .p0(node_level1_pos117_outp), .g0(node_level1_pos117_outg), .gp(node_level2_pos119_outg), .pp(node_level2_pos119_outp));
	wire node_level2_pos123_outg;
	wire node_level2_pos123_outp;
	pos_operator node_level2_pos123(.p1(node_level1_pos123_outp), .g1(node_level1_pos123_outg), .p0(node_level1_pos121_outp), .g0(node_level1_pos121_outg), .gp(node_level2_pos123_outg), .pp(node_level2_pos123_outp));
	wire node_level2_pos127_outg;
	wire node_level2_pos127_outp;
	pos_operator node_level2_pos127(.p1(node_level1_pos127_outp), .g1(node_level1_pos127_outg), .p0(node_level1_pos125_outp), .g0(node_level1_pos125_outg), .gp(node_level2_pos127_outg), .pp(node_level2_pos127_outp));
	wire node_level3_pos7_outg;
	wire node_level3_pos7_outp;
	neg_operator node_level3_pos7(.p1(node_level2_pos7_outp), .g1(node_level2_pos7_outg), .p0(node_level2_pos3_outp), .g0(node_level2_pos3_outg), .gp(node_level3_pos7_outg), .pp(node_level3_pos7_outp));
	wire node_level3_pos15_outg;
	wire node_level3_pos15_outp;
	neg_operator node_level3_pos15(.p1(node_level2_pos15_outp), .g1(node_level2_pos15_outg), .p0(node_level2_pos11_outp), .g0(node_level2_pos11_outg), .gp(node_level3_pos15_outg), .pp(node_level3_pos15_outp));
	wire node_level3_pos23_outg;
	wire node_level3_pos23_outp;
	neg_operator node_level3_pos23(.p1(node_level2_pos23_outp), .g1(node_level2_pos23_outg), .p0(node_level2_pos19_outp), .g0(node_level2_pos19_outg), .gp(node_level3_pos23_outg), .pp(node_level3_pos23_outp));
	wire node_level3_pos31_outg;
	wire node_level3_pos31_outp;
	neg_operator node_level3_pos31(.p1(node_level2_pos31_outp), .g1(node_level2_pos31_outg), .p0(node_level2_pos27_outp), .g0(node_level2_pos27_outg), .gp(node_level3_pos31_outg), .pp(node_level3_pos31_outp));
	wire node_level3_pos39_outg;
	wire node_level3_pos39_outp;
	neg_operator node_level3_pos39(.p1(node_level2_pos39_outp), .g1(node_level2_pos39_outg), .p0(node_level2_pos35_outp), .g0(node_level2_pos35_outg), .gp(node_level3_pos39_outg), .pp(node_level3_pos39_outp));
	wire node_level3_pos47_outg;
	wire node_level3_pos47_outp;
	neg_operator node_level3_pos47(.p1(node_level2_pos47_outp), .g1(node_level2_pos47_outg), .p0(node_level2_pos43_outp), .g0(node_level2_pos43_outg), .gp(node_level3_pos47_outg), .pp(node_level3_pos47_outp));
	wire node_level3_pos55_outg;
	wire node_level3_pos55_outp;
	neg_operator node_level3_pos55(.p1(node_level2_pos55_outp), .g1(node_level2_pos55_outg), .p0(node_level2_pos51_outp), .g0(node_level2_pos51_outg), .gp(node_level3_pos55_outg), .pp(node_level3_pos55_outp));
	wire node_level3_pos63_outg;
	wire node_level3_pos63_outp;
	neg_operator node_level3_pos63(.p1(node_level2_pos63_outp), .g1(node_level2_pos63_outg), .p0(node_level2_pos59_outp), .g0(node_level2_pos59_outg), .gp(node_level3_pos63_outg), .pp(node_level3_pos63_outp));
	wire node_level3_pos71_outg;
	wire node_level3_pos71_outp;
	neg_operator node_level3_pos71(.p1(node_level2_pos71_outp), .g1(node_level2_pos71_outg), .p0(node_level2_pos67_outp), .g0(node_level2_pos67_outg), .gp(node_level3_pos71_outg), .pp(node_level3_pos71_outp));
	wire node_level3_pos79_outg;
	wire node_level3_pos79_outp;
	neg_operator node_level3_pos79(.p1(node_level2_pos79_outp), .g1(node_level2_pos79_outg), .p0(node_level2_pos75_outp), .g0(node_level2_pos75_outg), .gp(node_level3_pos79_outg), .pp(node_level3_pos79_outp));
	wire node_level3_pos87_outg;
	wire node_level3_pos87_outp;
	neg_operator node_level3_pos87(.p1(node_level2_pos87_outp), .g1(node_level2_pos87_outg), .p0(node_level2_pos83_outp), .g0(node_level2_pos83_outg), .gp(node_level3_pos87_outg), .pp(node_level3_pos87_outp));
	wire node_level3_pos95_outg;
	wire node_level3_pos95_outp;
	neg_operator node_level3_pos95(.p1(node_level2_pos95_outp), .g1(node_level2_pos95_outg), .p0(node_level2_pos91_outp), .g0(node_level2_pos91_outg), .gp(node_level3_pos95_outg), .pp(node_level3_pos95_outp));
	wire node_level3_pos103_outg;
	wire node_level3_pos103_outp;
	neg_operator node_level3_pos103(.p1(node_level2_pos103_outp), .g1(node_level2_pos103_outg), .p0(node_level2_pos99_outp), .g0(node_level2_pos99_outg), .gp(node_level3_pos103_outg), .pp(node_level3_pos103_outp));
	wire node_level3_pos111_outg;
	wire node_level3_pos111_outp;
	neg_operator node_level3_pos111(.p1(node_level2_pos111_outp), .g1(node_level2_pos111_outg), .p0(node_level2_pos107_outp), .g0(node_level2_pos107_outg), .gp(node_level3_pos111_outg), .pp(node_level3_pos111_outp));
	wire node_level3_pos119_outg;
	wire node_level3_pos119_outp;
	neg_operator node_level3_pos119(.p1(node_level2_pos119_outp), .g1(node_level2_pos119_outg), .p0(node_level2_pos115_outp), .g0(node_level2_pos115_outg), .gp(node_level3_pos119_outg), .pp(node_level3_pos119_outp));
	wire node_level3_pos127_outg;
	wire node_level3_pos127_outp;
	neg_operator node_level3_pos127(.p1(node_level2_pos127_outp), .g1(node_level2_pos127_outg), .p0(node_level2_pos123_outp), .g0(node_level2_pos123_outg), .gp(node_level3_pos127_outg), .pp(node_level3_pos127_outp));
	wire node_level4_pos15_outg;
	wire node_level4_pos15_outp;
	pos_operator node_level4_pos15(.p1(node_level3_pos15_outp), .g1(node_level3_pos15_outg), .p0(node_level3_pos7_outp), .g0(node_level3_pos7_outg), .gp(node_level4_pos15_outg), .pp(node_level4_pos15_outp));
	wire node_level4_pos31_outg;
	wire node_level4_pos31_outp;
	pos_operator node_level4_pos31(.p1(node_level3_pos31_outp), .g1(node_level3_pos31_outg), .p0(node_level3_pos23_outp), .g0(node_level3_pos23_outg), .gp(node_level4_pos31_outg), .pp(node_level4_pos31_outp));
	wire node_level4_pos47_outg;
	wire node_level4_pos47_outp;
	pos_operator node_level4_pos47(.p1(node_level3_pos47_outp), .g1(node_level3_pos47_outg), .p0(node_level3_pos39_outp), .g0(node_level3_pos39_outg), .gp(node_level4_pos47_outg), .pp(node_level4_pos47_outp));
	wire node_level4_pos63_outg;
	wire node_level4_pos63_outp;
	pos_operator node_level4_pos63(.p1(node_level3_pos63_outp), .g1(node_level3_pos63_outg), .p0(node_level3_pos55_outp), .g0(node_level3_pos55_outg), .gp(node_level4_pos63_outg), .pp(node_level4_pos63_outp));
	wire node_level4_pos79_outg;
	wire node_level4_pos79_outp;
	pos_operator node_level4_pos79(.p1(node_level3_pos79_outp), .g1(node_level3_pos79_outg), .p0(node_level3_pos71_outp), .g0(node_level3_pos71_outg), .gp(node_level4_pos79_outg), .pp(node_level4_pos79_outp));
	wire node_level4_pos95_outg;
	wire node_level4_pos95_outp;
	pos_operator node_level4_pos95(.p1(node_level3_pos95_outp), .g1(node_level3_pos95_outg), .p0(node_level3_pos87_outp), .g0(node_level3_pos87_outg), .gp(node_level4_pos95_outg), .pp(node_level4_pos95_outp));
	wire node_level4_pos111_outg;
	wire node_level4_pos111_outp;
	pos_operator node_level4_pos111(.p1(node_level3_pos111_outp), .g1(node_level3_pos111_outg), .p0(node_level3_pos103_outp), .g0(node_level3_pos103_outg), .gp(node_level4_pos111_outg), .pp(node_level4_pos111_outp));
	wire node_level4_pos127_outg;
	wire node_level4_pos127_outp;
	pos_operator node_level4_pos127(.p1(node_level3_pos127_outp), .g1(node_level3_pos127_outg), .p0(node_level3_pos119_outp), .g0(node_level3_pos119_outg), .gp(node_level4_pos127_outg), .pp(node_level4_pos127_outp));
	wire node_level5_pos31_outg;
	wire node_level5_pos31_outp;
	neg_operator node_level5_pos31(.p1(node_level4_pos31_outp), .g1(node_level4_pos31_outg), .p0(node_level4_pos15_outp), .g0(node_level4_pos15_outg), .gp(node_level5_pos31_outg), .pp(node_level5_pos31_outp));
	wire node_level5_pos47_outg;
	wire node_level5_pos47_outp;
	neg_operator node_level5_pos47(.p1(node_level4_pos47_outp), .g1(node_level4_pos47_outg), .p0(node_level4_pos31_outp), .g0(node_level4_pos31_outg), .gp(node_level5_pos47_outg), .pp(node_level5_pos47_outp));
	wire node_level5_pos63_outg;
	wire node_level5_pos63_outp;
	neg_operator node_level5_pos63(.p1(node_level4_pos63_outp), .g1(node_level4_pos63_outg), .p0(node_level4_pos47_outp), .g0(node_level4_pos47_outg), .gp(node_level5_pos63_outg), .pp(node_level5_pos63_outp));
	wire node_level5_pos79_outg;
	wire node_level5_pos79_outp;
	neg_operator node_level5_pos79(.p1(node_level4_pos79_outp), .g1(node_level4_pos79_outg), .p0(node_level4_pos63_outp), .g0(node_level4_pos63_outg), .gp(node_level5_pos79_outg), .pp(node_level5_pos79_outp));
	wire node_level5_pos95_outg;
	wire node_level5_pos95_outp;
	neg_operator node_level5_pos95(.p1(node_level4_pos95_outp), .g1(node_level4_pos95_outg), .p0(node_level4_pos79_outp), .g0(node_level4_pos79_outg), .gp(node_level5_pos95_outg), .pp(node_level5_pos95_outp));
	wire node_level5_pos111_outg;
	wire node_level5_pos111_outp;
	neg_operator node_level5_pos111(.p1(node_level4_pos111_outp), .g1(node_level4_pos111_outg), .p0(node_level4_pos95_outp), .g0(node_level4_pos95_outg), .gp(node_level5_pos111_outg), .pp(node_level5_pos111_outp));
	wire node_level5_pos127_outg;
	wire node_level5_pos127_outp;
	neg_operator node_level5_pos127(.p1(node_level4_pos127_outp), .g1(node_level4_pos127_outg), .p0(node_level4_pos111_outp), .g0(node_level4_pos111_outg), .gp(node_level5_pos127_outg), .pp(node_level5_pos127_outp));
	wire node_level6_pos47_outg;
	wire node_level6_pos47_outp;
	pos_operator node_level6_pos47(.p1(node_level5_pos47_outp), .g1(node_level5_pos47_outg), .p0(~node_level4_pos15_outp), .g0(~node_level4_pos15_outg), .gp(node_level6_pos47_outg), .pp(node_level6_pos47_outp));
	wire node_level6_pos63_outg;
	wire node_level6_pos63_outp;
	pos_operator node_level6_pos63(.p1(node_level5_pos63_outp), .g1(node_level5_pos63_outg), .p0(node_level5_pos31_outp), .g0(node_level5_pos31_outg), .gp(node_level6_pos63_outg), .pp(node_level6_pos63_outp));
	wire node_level6_pos79_outg;
	wire node_level6_pos79_outp;
	pos_operator node_level6_pos79(.p1(node_level5_pos79_outp), .g1(node_level5_pos79_outg), .p0(node_level5_pos47_outp), .g0(node_level5_pos47_outg), .gp(node_level6_pos79_outg), .pp(node_level6_pos79_outp));
	wire node_level6_pos95_outg;
	wire node_level6_pos95_outp;
	pos_operator node_level6_pos95(.p1(node_level5_pos95_outp), .g1(node_level5_pos95_outg), .p0(node_level5_pos63_outp), .g0(node_level5_pos63_outg), .gp(node_level6_pos95_outg), .pp(node_level6_pos95_outp));
	wire node_level6_pos111_outg;
	wire node_level6_pos111_outp;
	pos_operator node_level6_pos111(.p1(node_level5_pos111_outp), .g1(node_level5_pos111_outg), .p0(node_level5_pos79_outp), .g0(node_level5_pos79_outg), .gp(node_level6_pos111_outg), .pp(node_level6_pos111_outp));
	wire node_level6_pos127_outg;
	wire node_level6_pos127_outp;
	pos_operator node_level6_pos127(.p1(node_level5_pos127_outp), .g1(node_level5_pos127_outg), .p0(node_level5_pos95_outp), .g0(node_level5_pos95_outg), .gp(node_level6_pos127_outg), .pp(node_level6_pos127_outp));
	wire node_level7_pos79_outg;
	wire node_level7_pos79_outp;
	neg_operator node_level7_pos79(.p1(node_level6_pos79_outp), .g1(node_level6_pos79_outg), .p0(node_level4_pos15_outp), .g0(node_level4_pos15_outg), .gp(node_level7_pos79_outg), .pp(node_level7_pos79_outp));
	wire node_level7_pos95_outg;
	wire node_level7_pos95_outp;
	neg_operator node_level7_pos95(.p1(node_level6_pos95_outp), .g1(node_level6_pos95_outg), .p0(~node_level5_pos31_outp), .g0(~node_level5_pos31_outg), .gp(node_level7_pos95_outg), .pp(node_level7_pos95_outp));
	wire node_level7_pos111_outg;
	wire node_level7_pos111_outp;
	neg_operator node_level7_pos111(.p1(node_level6_pos111_outp), .g1(node_level6_pos111_outg), .p0(node_level6_pos47_outp), .g0(node_level6_pos47_outg), .gp(node_level7_pos111_outg), .pp(node_level7_pos111_outp));
	wire node_level7_pos127_outg;
	wire node_level7_pos127_outp;
	neg_operator node_level7_pos127(.p1(node_level6_pos127_outp), .g1(node_level6_pos127_outg), .p0(node_level6_pos63_outp), .g0(node_level6_pos63_outg), .gp(node_level7_pos127_outg), .pp(node_level7_pos127_outp));
	wire node_level8_pos23_outg;
	wire node_level8_pos23_outp;
	pos_operator node_level8_pos23(.p1(node_level3_pos23_outp), .g1(node_level3_pos23_outg), .p0(~node_level4_pos15_outp), .g0(~node_level4_pos15_outg), .gp(node_level8_pos23_outg), .pp(node_level8_pos23_outp));
	wire node_level8_pos39_outg;
	wire node_level8_pos39_outp;
	pos_operator node_level8_pos39(.p1(node_level3_pos39_outp), .g1(node_level3_pos39_outg), .p0(node_level5_pos31_outp), .g0(node_level5_pos31_outg), .gp(node_level8_pos39_outg), .pp(node_level8_pos39_outp));
	wire node_level8_pos55_outg;
	wire node_level8_pos55_outp;
	pos_operator node_level8_pos55(.p1(node_level3_pos55_outp), .g1(node_level3_pos55_outg), .p0(~node_level6_pos47_outp), .g0(~node_level6_pos47_outg), .gp(node_level8_pos55_outg), .pp(node_level8_pos55_outp));
	wire node_level8_pos71_outg;
	wire node_level8_pos71_outp;
	pos_operator node_level8_pos71(.p1(node_level3_pos71_outp), .g1(node_level3_pos71_outg), .p0(~node_level6_pos63_outp), .g0(~node_level6_pos63_outg), .gp(node_level8_pos71_outg), .pp(node_level8_pos71_outp));
	wire node_level8_pos87_outg;
	wire node_level8_pos87_outp;
	pos_operator node_level8_pos87(.p1(node_level3_pos87_outp), .g1(node_level3_pos87_outg), .p0(node_level7_pos79_outp), .g0(node_level7_pos79_outg), .gp(node_level8_pos87_outg), .pp(node_level8_pos87_outp));
	wire node_level8_pos103_outg;
	wire node_level8_pos103_outp;
	pos_operator node_level8_pos103(.p1(node_level3_pos103_outp), .g1(node_level3_pos103_outg), .p0(node_level7_pos95_outp), .g0(node_level7_pos95_outg), .gp(node_level8_pos103_outg), .pp(node_level8_pos103_outp));
	wire node_level8_pos119_outg;
	wire node_level8_pos119_outp;
	pos_operator node_level8_pos119(.p1(node_level3_pos119_outp), .g1(node_level3_pos119_outg), .p0(node_level7_pos111_outp), .g0(node_level7_pos111_outg), .gp(node_level8_pos119_outg), .pp(node_level8_pos119_outp));
	wire node_level9_pos11_outg;
	wire node_level9_pos11_outp;
	neg_operator node_level9_pos11(.p1(node_level2_pos11_outp), .g1(node_level2_pos11_outg), .p0(~node_level3_pos7_outp), .g0(~node_level3_pos7_outg), .gp(node_level9_pos11_outg), .pp(node_level9_pos11_outp));
	wire node_level9_pos19_outg;
	wire node_level9_pos19_outp;
	neg_operator node_level9_pos19(.p1(node_level2_pos19_outp), .g1(node_level2_pos19_outg), .p0(node_level4_pos15_outp), .g0(node_level4_pos15_outg), .gp(node_level9_pos19_outg), .pp(node_level9_pos19_outp));
	wire node_level9_pos27_outg;
	wire node_level9_pos27_outp;
	neg_operator node_level9_pos27(.p1(node_level2_pos27_outp), .g1(node_level2_pos27_outg), .p0(node_level8_pos23_outp), .g0(node_level8_pos23_outg), .gp(node_level9_pos27_outg), .pp(node_level9_pos27_outp));
	wire node_level9_pos35_outg;
	wire node_level9_pos35_outp;
	neg_operator node_level9_pos35(.p1(node_level2_pos35_outp), .g1(node_level2_pos35_outg), .p0(~node_level5_pos31_outp), .g0(~node_level5_pos31_outg), .gp(node_level9_pos35_outg), .pp(node_level9_pos35_outp));
	wire node_level9_pos43_outg;
	wire node_level9_pos43_outp;
	neg_operator node_level9_pos43(.p1(node_level2_pos43_outp), .g1(node_level2_pos43_outg), .p0(node_level8_pos39_outp), .g0(node_level8_pos39_outg), .gp(node_level9_pos43_outg), .pp(node_level9_pos43_outp));
	wire node_level9_pos51_outg;
	wire node_level9_pos51_outp;
	neg_operator node_level9_pos51(.p1(node_level2_pos51_outp), .g1(node_level2_pos51_outg), .p0(node_level6_pos47_outp), .g0(node_level6_pos47_outg), .gp(node_level9_pos51_outg), .pp(node_level9_pos51_outp));
	wire node_level9_pos59_outg;
	wire node_level9_pos59_outp;
	neg_operator node_level9_pos59(.p1(node_level2_pos59_outp), .g1(node_level2_pos59_outg), .p0(node_level8_pos55_outp), .g0(node_level8_pos55_outg), .gp(node_level9_pos59_outg), .pp(node_level9_pos59_outp));
	wire node_level9_pos67_outg;
	wire node_level9_pos67_outp;
	neg_operator node_level9_pos67(.p1(node_level2_pos67_outp), .g1(node_level2_pos67_outg), .p0(node_level6_pos63_outp), .g0(node_level6_pos63_outg), .gp(node_level9_pos67_outg), .pp(node_level9_pos67_outp));
	wire node_level9_pos75_outg;
	wire node_level9_pos75_outp;
	neg_operator node_level9_pos75(.p1(node_level2_pos75_outp), .g1(node_level2_pos75_outg), .p0(node_level8_pos71_outp), .g0(node_level8_pos71_outg), .gp(node_level9_pos75_outg), .pp(node_level9_pos75_outp));
	wire node_level9_pos83_outg;
	wire node_level9_pos83_outp;
	neg_operator node_level9_pos83(.p1(node_level2_pos83_outp), .g1(node_level2_pos83_outg), .p0(~node_level7_pos79_outp), .g0(~node_level7_pos79_outg), .gp(node_level9_pos83_outg), .pp(node_level9_pos83_outp));
	wire node_level9_pos91_outg;
	wire node_level9_pos91_outp;
	neg_operator node_level9_pos91(.p1(node_level2_pos91_outp), .g1(node_level2_pos91_outg), .p0(node_level8_pos87_outp), .g0(node_level8_pos87_outg), .gp(node_level9_pos91_outg), .pp(node_level9_pos91_outp));
	wire node_level9_pos99_outg;
	wire node_level9_pos99_outp;
	neg_operator node_level9_pos99(.p1(node_level2_pos99_outp), .g1(node_level2_pos99_outg), .p0(~node_level7_pos95_outp), .g0(~node_level7_pos95_outg), .gp(node_level9_pos99_outg), .pp(node_level9_pos99_outp));
	wire node_level9_pos107_outg;
	wire node_level9_pos107_outp;
	neg_operator node_level9_pos107(.p1(node_level2_pos107_outp), .g1(node_level2_pos107_outg), .p0(node_level8_pos103_outp), .g0(node_level8_pos103_outg), .gp(node_level9_pos107_outg), .pp(node_level9_pos107_outp));
	wire node_level9_pos115_outg;
	wire node_level9_pos115_outp;
	neg_operator node_level9_pos115(.p1(node_level2_pos115_outp), .g1(node_level2_pos115_outg), .p0(~node_level7_pos111_outp), .g0(~node_level7_pos111_outg), .gp(node_level9_pos115_outg), .pp(node_level9_pos115_outp));
	wire node_level9_pos123_outg;
	wire node_level9_pos123_outp;
	neg_operator node_level9_pos123(.p1(node_level2_pos123_outp), .g1(node_level2_pos123_outg), .p0(node_level8_pos119_outp), .g0(node_level8_pos119_outg), .gp(node_level9_pos123_outg), .pp(node_level9_pos123_outp));
	wire node_level10_pos5_outg;
	wire node_level10_pos5_outp;
	pos_operator node_level10_pos5(.p1(node_level1_pos5_outp), .g1(node_level1_pos5_outg), .p0(~node_level2_pos3_outp), .g0(~node_level2_pos3_outg), .gp(node_level10_pos5_outg), .pp(node_level10_pos5_outp));
	wire node_level10_pos9_outg;
	wire node_level10_pos9_outp;
	pos_operator node_level10_pos9(.p1(node_level1_pos9_outp), .g1(node_level1_pos9_outg), .p0(node_level3_pos7_outp), .g0(node_level3_pos7_outg), .gp(node_level10_pos9_outg), .pp(node_level10_pos9_outp));
	wire node_level10_pos13_outg;
	wire node_level10_pos13_outp;
	pos_operator node_level10_pos13(.p1(node_level1_pos13_outp), .g1(node_level1_pos13_outg), .p0(node_level9_pos11_outp), .g0(node_level9_pos11_outg), .gp(node_level10_pos13_outg), .pp(node_level10_pos13_outp));
	wire node_level10_pos17_outg;
	wire node_level10_pos17_outp;
	pos_operator node_level10_pos17(.p1(node_level1_pos17_outp), .g1(node_level1_pos17_outg), .p0(~node_level4_pos15_outp), .g0(~node_level4_pos15_outg), .gp(node_level10_pos17_outg), .pp(node_level10_pos17_outp));
	wire node_level10_pos21_outg;
	wire node_level10_pos21_outp;
	pos_operator node_level10_pos21(.p1(node_level1_pos21_outp), .g1(node_level1_pos21_outg), .p0(node_level9_pos19_outp), .g0(node_level9_pos19_outg), .gp(node_level10_pos21_outg), .pp(node_level10_pos21_outp));
	wire node_level10_pos25_outg;
	wire node_level10_pos25_outp;
	pos_operator node_level10_pos25(.p1(node_level1_pos25_outp), .g1(node_level1_pos25_outg), .p0(~node_level8_pos23_outp), .g0(~node_level8_pos23_outg), .gp(node_level10_pos25_outg), .pp(node_level10_pos25_outp));
	wire node_level10_pos29_outg;
	wire node_level10_pos29_outp;
	pos_operator node_level10_pos29(.p1(node_level1_pos29_outp), .g1(node_level1_pos29_outg), .p0(node_level9_pos27_outp), .g0(node_level9_pos27_outg), .gp(node_level10_pos29_outg), .pp(node_level10_pos29_outp));
	wire node_level10_pos33_outg;
	wire node_level10_pos33_outp;
	pos_operator node_level10_pos33(.p1(node_level1_pos33_outp), .g1(node_level1_pos33_outg), .p0(node_level5_pos31_outp), .g0(node_level5_pos31_outg), .gp(node_level10_pos33_outg), .pp(node_level10_pos33_outp));
	wire node_level10_pos37_outg;
	wire node_level10_pos37_outp;
	pos_operator node_level10_pos37(.p1(node_level1_pos37_outp), .g1(node_level1_pos37_outg), .p0(node_level9_pos35_outp), .g0(node_level9_pos35_outg), .gp(node_level10_pos37_outg), .pp(node_level10_pos37_outp));
	wire node_level10_pos41_outg;
	wire node_level10_pos41_outp;
	pos_operator node_level10_pos41(.p1(node_level1_pos41_outp), .g1(node_level1_pos41_outg), .p0(~node_level8_pos39_outp), .g0(~node_level8_pos39_outg), .gp(node_level10_pos41_outg), .pp(node_level10_pos41_outp));
	wire node_level10_pos45_outg;
	wire node_level10_pos45_outp;
	pos_operator node_level10_pos45(.p1(node_level1_pos45_outp), .g1(node_level1_pos45_outg), .p0(node_level9_pos43_outp), .g0(node_level9_pos43_outg), .gp(node_level10_pos45_outg), .pp(node_level10_pos45_outp));
	wire node_level10_pos49_outg;
	wire node_level10_pos49_outp;
	pos_operator node_level10_pos49(.p1(node_level1_pos49_outp), .g1(node_level1_pos49_outg), .p0(~node_level6_pos47_outp), .g0(~node_level6_pos47_outg), .gp(node_level10_pos49_outg), .pp(node_level10_pos49_outp));
	wire node_level10_pos53_outg;
	wire node_level10_pos53_outp;
	pos_operator node_level10_pos53(.p1(node_level1_pos53_outp), .g1(node_level1_pos53_outg), .p0(node_level9_pos51_outp), .g0(node_level9_pos51_outg), .gp(node_level10_pos53_outg), .pp(node_level10_pos53_outp));
	wire node_level10_pos57_outg;
	wire node_level10_pos57_outp;
	pos_operator node_level10_pos57(.p1(node_level1_pos57_outp), .g1(node_level1_pos57_outg), .p0(~node_level8_pos55_outp), .g0(~node_level8_pos55_outg), .gp(node_level10_pos57_outg), .pp(node_level10_pos57_outp));
	wire node_level10_pos61_outg;
	wire node_level10_pos61_outp;
	pos_operator node_level10_pos61(.p1(node_level1_pos61_outp), .g1(node_level1_pos61_outg), .p0(node_level9_pos59_outp), .g0(node_level9_pos59_outg), .gp(node_level10_pos61_outg), .pp(node_level10_pos61_outp));
	wire node_level10_pos65_outg;
	wire node_level10_pos65_outp;
	pos_operator node_level10_pos65(.p1(node_level1_pos65_outp), .g1(node_level1_pos65_outg), .p0(~node_level6_pos63_outp), .g0(~node_level6_pos63_outg), .gp(node_level10_pos65_outg), .pp(node_level10_pos65_outp));
	wire node_level10_pos69_outg;
	wire node_level10_pos69_outp;
	pos_operator node_level10_pos69(.p1(node_level1_pos69_outp), .g1(node_level1_pos69_outg), .p0(node_level9_pos67_outp), .g0(node_level9_pos67_outg), .gp(node_level10_pos69_outg), .pp(node_level10_pos69_outp));
	wire node_level10_pos73_outg;
	wire node_level10_pos73_outp;
	pos_operator node_level10_pos73(.p1(node_level1_pos73_outp), .g1(node_level1_pos73_outg), .p0(~node_level8_pos71_outp), .g0(~node_level8_pos71_outg), .gp(node_level10_pos73_outg), .pp(node_level10_pos73_outp));
	wire node_level10_pos77_outg;
	wire node_level10_pos77_outp;
	pos_operator node_level10_pos77(.p1(node_level1_pos77_outp), .g1(node_level1_pos77_outg), .p0(node_level9_pos75_outp), .g0(node_level9_pos75_outg), .gp(node_level10_pos77_outg), .pp(node_level10_pos77_outp));
	wire node_level10_pos81_outg;
	wire node_level10_pos81_outp;
	pos_operator node_level10_pos81(.p1(node_level1_pos81_outp), .g1(node_level1_pos81_outg), .p0(node_level7_pos79_outp), .g0(node_level7_pos79_outg), .gp(node_level10_pos81_outg), .pp(node_level10_pos81_outp));
	wire node_level10_pos85_outg;
	wire node_level10_pos85_outp;
	pos_operator node_level10_pos85(.p1(node_level1_pos85_outp), .g1(node_level1_pos85_outg), .p0(node_level9_pos83_outp), .g0(node_level9_pos83_outg), .gp(node_level10_pos85_outg), .pp(node_level10_pos85_outp));
	wire node_level10_pos89_outg;
	wire node_level10_pos89_outp;
	pos_operator node_level10_pos89(.p1(node_level1_pos89_outp), .g1(node_level1_pos89_outg), .p0(~node_level8_pos87_outp), .g0(~node_level8_pos87_outg), .gp(node_level10_pos89_outg), .pp(node_level10_pos89_outp));
	wire node_level10_pos93_outg;
	wire node_level10_pos93_outp;
	pos_operator node_level10_pos93(.p1(node_level1_pos93_outp), .g1(node_level1_pos93_outg), .p0(node_level9_pos91_outp), .g0(node_level9_pos91_outg), .gp(node_level10_pos93_outg), .pp(node_level10_pos93_outp));
	wire node_level10_pos97_outg;
	wire node_level10_pos97_outp;
	pos_operator node_level10_pos97(.p1(node_level1_pos97_outp), .g1(node_level1_pos97_outg), .p0(node_level7_pos95_outp), .g0(node_level7_pos95_outg), .gp(node_level10_pos97_outg), .pp(node_level10_pos97_outp));
	wire node_level10_pos101_outg;
	wire node_level10_pos101_outp;
	pos_operator node_level10_pos101(.p1(node_level1_pos101_outp), .g1(node_level1_pos101_outg), .p0(node_level9_pos99_outp), .g0(node_level9_pos99_outg), .gp(node_level10_pos101_outg), .pp(node_level10_pos101_outp));
	wire node_level10_pos105_outg;
	wire node_level10_pos105_outp;
	pos_operator node_level10_pos105(.p1(node_level1_pos105_outp), .g1(node_level1_pos105_outg), .p0(~node_level8_pos103_outp), .g0(~node_level8_pos103_outg), .gp(node_level10_pos105_outg), .pp(node_level10_pos105_outp));
	wire node_level10_pos109_outg;
	wire node_level10_pos109_outp;
	pos_operator node_level10_pos109(.p1(node_level1_pos109_outp), .g1(node_level1_pos109_outg), .p0(node_level9_pos107_outp), .g0(node_level9_pos107_outg), .gp(node_level10_pos109_outg), .pp(node_level10_pos109_outp));
	wire node_level10_pos113_outg;
	wire node_level10_pos113_outp;
	pos_operator node_level10_pos113(.p1(node_level1_pos113_outp), .g1(node_level1_pos113_outg), .p0(node_level7_pos111_outp), .g0(node_level7_pos111_outg), .gp(node_level10_pos113_outg), .pp(node_level10_pos113_outp));
	wire node_level10_pos117_outg;
	wire node_level10_pos117_outp;
	pos_operator node_level10_pos117(.p1(node_level1_pos117_outp), .g1(node_level1_pos117_outg), .p0(node_level9_pos115_outp), .g0(node_level9_pos115_outg), .gp(node_level10_pos117_outg), .pp(node_level10_pos117_outp));
	wire node_level10_pos121_outg;
	wire node_level10_pos121_outp;
	pos_operator node_level10_pos121(.p1(node_level1_pos121_outp), .g1(node_level1_pos121_outg), .p0(~node_level8_pos119_outp), .g0(~node_level8_pos119_outg), .gp(node_level10_pos121_outg), .pp(node_level10_pos121_outp));
	wire node_level10_pos125_outg;
	wire node_level10_pos125_outp;
	pos_operator node_level10_pos125(.p1(node_level1_pos125_outp), .g1(node_level1_pos125_outg), .p0(node_level9_pos123_outp), .g0(node_level9_pos123_outg), .gp(node_level10_pos125_outg), .pp(node_level10_pos125_outp));
	wire node_level11_pos2_outg;
	wire node_level11_pos2_outp;
	neg_operator node_level11_pos2(.p1(p_in[2]), .g1(g_in[2]), .p0(~node_level1_pos1_outp), .g0(~node_level1_pos1_outg), .gp(node_level11_pos2_outg), .pp(node_level11_pos2_outp));
	wire node_level11_pos4_outg;
	wire node_level11_pos4_outp;
	neg_operator node_level11_pos4(.p1(p_in[4]), .g1(g_in[4]), .p0(node_level2_pos3_outp), .g0(node_level2_pos3_outg), .gp(node_level11_pos4_outg), .pp(node_level11_pos4_outp));
	wire node_level11_pos6_outg;
	wire node_level11_pos6_outp;
	neg_operator node_level11_pos6(.p1(p_in[6]), .g1(g_in[6]), .p0(node_level10_pos5_outp), .g0(node_level10_pos5_outg), .gp(node_level11_pos6_outg), .pp(node_level11_pos6_outp));
	wire node_level11_pos8_outg;
	wire node_level11_pos8_outp;
	neg_operator node_level11_pos8(.p1(p_in[8]), .g1(g_in[8]), .p0(~node_level3_pos7_outp), .g0(~node_level3_pos7_outg), .gp(node_level11_pos8_outg), .pp(node_level11_pos8_outp));
	wire node_level11_pos10_outg;
	wire node_level11_pos10_outp;
	neg_operator node_level11_pos10(.p1(p_in[10]), .g1(g_in[10]), .p0(node_level10_pos9_outp), .g0(node_level10_pos9_outg), .gp(node_level11_pos10_outg), .pp(node_level11_pos10_outp));
	wire node_level11_pos12_outg;
	wire node_level11_pos12_outp;
	neg_operator node_level11_pos12(.p1(p_in[12]), .g1(g_in[12]), .p0(~node_level9_pos11_outp), .g0(~node_level9_pos11_outg), .gp(node_level11_pos12_outg), .pp(node_level11_pos12_outp));
	wire node_level11_pos14_outg;
	wire node_level11_pos14_outp;
	neg_operator node_level11_pos14(.p1(p_in[14]), .g1(g_in[14]), .p0(node_level10_pos13_outp), .g0(node_level10_pos13_outg), .gp(node_level11_pos14_outg), .pp(node_level11_pos14_outp));
	wire node_level11_pos16_outg;
	wire node_level11_pos16_outp;
	neg_operator node_level11_pos16(.p1(p_in[16]), .g1(g_in[16]), .p0(node_level4_pos15_outp), .g0(node_level4_pos15_outg), .gp(node_level11_pos16_outg), .pp(node_level11_pos16_outp));
	wire node_level11_pos18_outg;
	wire node_level11_pos18_outp;
	neg_operator node_level11_pos18(.p1(p_in[18]), .g1(g_in[18]), .p0(node_level10_pos17_outp), .g0(node_level10_pos17_outg), .gp(node_level11_pos18_outg), .pp(node_level11_pos18_outp));
	wire node_level11_pos20_outg;
	wire node_level11_pos20_outp;
	neg_operator node_level11_pos20(.p1(p_in[20]), .g1(g_in[20]), .p0(~node_level9_pos19_outp), .g0(~node_level9_pos19_outg), .gp(node_level11_pos20_outg), .pp(node_level11_pos20_outp));
	wire node_level11_pos22_outg;
	wire node_level11_pos22_outp;
	neg_operator node_level11_pos22(.p1(p_in[22]), .g1(g_in[22]), .p0(node_level10_pos21_outp), .g0(node_level10_pos21_outg), .gp(node_level11_pos22_outg), .pp(node_level11_pos22_outp));
	wire node_level11_pos24_outg;
	wire node_level11_pos24_outp;
	neg_operator node_level11_pos24(.p1(p_in[24]), .g1(g_in[24]), .p0(node_level8_pos23_outp), .g0(node_level8_pos23_outg), .gp(node_level11_pos24_outg), .pp(node_level11_pos24_outp));
	wire node_level11_pos26_outg;
	wire node_level11_pos26_outp;
	neg_operator node_level11_pos26(.p1(p_in[26]), .g1(g_in[26]), .p0(node_level10_pos25_outp), .g0(node_level10_pos25_outg), .gp(node_level11_pos26_outg), .pp(node_level11_pos26_outp));
	wire node_level11_pos28_outg;
	wire node_level11_pos28_outp;
	neg_operator node_level11_pos28(.p1(p_in[28]), .g1(g_in[28]), .p0(~node_level9_pos27_outp), .g0(~node_level9_pos27_outg), .gp(node_level11_pos28_outg), .pp(node_level11_pos28_outp));
	wire node_level11_pos30_outg;
	wire node_level11_pos30_outp;
	neg_operator node_level11_pos30(.p1(p_in[30]), .g1(g_in[30]), .p0(node_level10_pos29_outp), .g0(node_level10_pos29_outg), .gp(node_level11_pos30_outg), .pp(node_level11_pos30_outp));
	wire node_level11_pos32_outg;
	wire node_level11_pos32_outp;
	neg_operator node_level11_pos32(.p1(p_in[32]), .g1(g_in[32]), .p0(~node_level5_pos31_outp), .g0(~node_level5_pos31_outg), .gp(node_level11_pos32_outg), .pp(node_level11_pos32_outp));
	wire node_level11_pos34_outg;
	wire node_level11_pos34_outp;
	neg_operator node_level11_pos34(.p1(p_in[34]), .g1(g_in[34]), .p0(node_level10_pos33_outp), .g0(node_level10_pos33_outg), .gp(node_level11_pos34_outg), .pp(node_level11_pos34_outp));
	wire node_level11_pos36_outg;
	wire node_level11_pos36_outp;
	neg_operator node_level11_pos36(.p1(p_in[36]), .g1(g_in[36]), .p0(~node_level9_pos35_outp), .g0(~node_level9_pos35_outg), .gp(node_level11_pos36_outg), .pp(node_level11_pos36_outp));
	wire node_level11_pos38_outg;
	wire node_level11_pos38_outp;
	neg_operator node_level11_pos38(.p1(p_in[38]), .g1(g_in[38]), .p0(node_level10_pos37_outp), .g0(node_level10_pos37_outg), .gp(node_level11_pos38_outg), .pp(node_level11_pos38_outp));
	wire node_level11_pos40_outg;
	wire node_level11_pos40_outp;
	neg_operator node_level11_pos40(.p1(p_in[40]), .g1(g_in[40]), .p0(node_level8_pos39_outp), .g0(node_level8_pos39_outg), .gp(node_level11_pos40_outg), .pp(node_level11_pos40_outp));
	wire node_level11_pos42_outg;
	wire node_level11_pos42_outp;
	neg_operator node_level11_pos42(.p1(p_in[42]), .g1(g_in[42]), .p0(node_level10_pos41_outp), .g0(node_level10_pos41_outg), .gp(node_level11_pos42_outg), .pp(node_level11_pos42_outp));
	wire node_level11_pos44_outg;
	wire node_level11_pos44_outp;
	neg_operator node_level11_pos44(.p1(p_in[44]), .g1(g_in[44]), .p0(~node_level9_pos43_outp), .g0(~node_level9_pos43_outg), .gp(node_level11_pos44_outg), .pp(node_level11_pos44_outp));
	wire node_level11_pos46_outg;
	wire node_level11_pos46_outp;
	neg_operator node_level11_pos46(.p1(p_in[46]), .g1(g_in[46]), .p0(node_level10_pos45_outp), .g0(node_level10_pos45_outg), .gp(node_level11_pos46_outg), .pp(node_level11_pos46_outp));
	wire node_level11_pos48_outg;
	wire node_level11_pos48_outp;
	neg_operator node_level11_pos48(.p1(p_in[48]), .g1(g_in[48]), .p0(node_level6_pos47_outp), .g0(node_level6_pos47_outg), .gp(node_level11_pos48_outg), .pp(node_level11_pos48_outp));
	wire node_level11_pos50_outg;
	wire node_level11_pos50_outp;
	neg_operator node_level11_pos50(.p1(p_in[50]), .g1(g_in[50]), .p0(node_level10_pos49_outp), .g0(node_level10_pos49_outg), .gp(node_level11_pos50_outg), .pp(node_level11_pos50_outp));
	wire node_level11_pos52_outg;
	wire node_level11_pos52_outp;
	neg_operator node_level11_pos52(.p1(p_in[52]), .g1(g_in[52]), .p0(~node_level9_pos51_outp), .g0(~node_level9_pos51_outg), .gp(node_level11_pos52_outg), .pp(node_level11_pos52_outp));
	wire node_level11_pos54_outg;
	wire node_level11_pos54_outp;
	neg_operator node_level11_pos54(.p1(p_in[54]), .g1(g_in[54]), .p0(node_level10_pos53_outp), .g0(node_level10_pos53_outg), .gp(node_level11_pos54_outg), .pp(node_level11_pos54_outp));
	wire node_level11_pos56_outg;
	wire node_level11_pos56_outp;
	neg_operator node_level11_pos56(.p1(p_in[56]), .g1(g_in[56]), .p0(node_level8_pos55_outp), .g0(node_level8_pos55_outg), .gp(node_level11_pos56_outg), .pp(node_level11_pos56_outp));
	wire node_level11_pos58_outg;
	wire node_level11_pos58_outp;
	neg_operator node_level11_pos58(.p1(p_in[58]), .g1(g_in[58]), .p0(node_level10_pos57_outp), .g0(node_level10_pos57_outg), .gp(node_level11_pos58_outg), .pp(node_level11_pos58_outp));
	wire node_level11_pos60_outg;
	wire node_level11_pos60_outp;
	neg_operator node_level11_pos60(.p1(p_in[60]), .g1(g_in[60]), .p0(~node_level9_pos59_outp), .g0(~node_level9_pos59_outg), .gp(node_level11_pos60_outg), .pp(node_level11_pos60_outp));
	wire node_level11_pos62_outg;
	wire node_level11_pos62_outp;
	neg_operator node_level11_pos62(.p1(p_in[62]), .g1(g_in[62]), .p0(node_level10_pos61_outp), .g0(node_level10_pos61_outg), .gp(node_level11_pos62_outg), .pp(node_level11_pos62_outp));
	wire node_level11_pos64_outg;
	wire node_level11_pos64_outp;
	neg_operator node_level11_pos64(.p1(p_in[64]), .g1(g_in[64]), .p0(node_level6_pos63_outp), .g0(node_level6_pos63_outg), .gp(node_level11_pos64_outg), .pp(node_level11_pos64_outp));
	wire node_level11_pos66_outg;
	wire node_level11_pos66_outp;
	neg_operator node_level11_pos66(.p1(p_in[66]), .g1(g_in[66]), .p0(node_level10_pos65_outp), .g0(node_level10_pos65_outg), .gp(node_level11_pos66_outg), .pp(node_level11_pos66_outp));
	wire node_level11_pos68_outg;
	wire node_level11_pos68_outp;
	neg_operator node_level11_pos68(.p1(p_in[68]), .g1(g_in[68]), .p0(~node_level9_pos67_outp), .g0(~node_level9_pos67_outg), .gp(node_level11_pos68_outg), .pp(node_level11_pos68_outp));
	wire node_level11_pos70_outg;
	wire node_level11_pos70_outp;
	neg_operator node_level11_pos70(.p1(p_in[70]), .g1(g_in[70]), .p0(node_level10_pos69_outp), .g0(node_level10_pos69_outg), .gp(node_level11_pos70_outg), .pp(node_level11_pos70_outp));
	wire node_level11_pos72_outg;
	wire node_level11_pos72_outp;
	neg_operator node_level11_pos72(.p1(p_in[72]), .g1(g_in[72]), .p0(node_level8_pos71_outp), .g0(node_level8_pos71_outg), .gp(node_level11_pos72_outg), .pp(node_level11_pos72_outp));
	wire node_level11_pos74_outg;
	wire node_level11_pos74_outp;
	neg_operator node_level11_pos74(.p1(p_in[74]), .g1(g_in[74]), .p0(node_level10_pos73_outp), .g0(node_level10_pos73_outg), .gp(node_level11_pos74_outg), .pp(node_level11_pos74_outp));
	wire node_level11_pos76_outg;
	wire node_level11_pos76_outp;
	neg_operator node_level11_pos76(.p1(p_in[76]), .g1(g_in[76]), .p0(~node_level9_pos75_outp), .g0(~node_level9_pos75_outg), .gp(node_level11_pos76_outg), .pp(node_level11_pos76_outp));
	wire node_level11_pos78_outg;
	wire node_level11_pos78_outp;
	neg_operator node_level11_pos78(.p1(p_in[78]), .g1(g_in[78]), .p0(node_level10_pos77_outp), .g0(node_level10_pos77_outg), .gp(node_level11_pos78_outg), .pp(node_level11_pos78_outp));
	wire node_level11_pos80_outg;
	wire node_level11_pos80_outp;
	neg_operator node_level11_pos80(.p1(p_in[80]), .g1(g_in[80]), .p0(~node_level7_pos79_outp), .g0(~node_level7_pos79_outg), .gp(node_level11_pos80_outg), .pp(node_level11_pos80_outp));
	wire node_level11_pos82_outg;
	wire node_level11_pos82_outp;
	neg_operator node_level11_pos82(.p1(p_in[82]), .g1(g_in[82]), .p0(node_level10_pos81_outp), .g0(node_level10_pos81_outg), .gp(node_level11_pos82_outg), .pp(node_level11_pos82_outp));
	wire node_level11_pos84_outg;
	wire node_level11_pos84_outp;
	neg_operator node_level11_pos84(.p1(p_in[84]), .g1(g_in[84]), .p0(~node_level9_pos83_outp), .g0(~node_level9_pos83_outg), .gp(node_level11_pos84_outg), .pp(node_level11_pos84_outp));
	wire node_level11_pos86_outg;
	wire node_level11_pos86_outp;
	neg_operator node_level11_pos86(.p1(p_in[86]), .g1(g_in[86]), .p0(node_level10_pos85_outp), .g0(node_level10_pos85_outg), .gp(node_level11_pos86_outg), .pp(node_level11_pos86_outp));
	wire node_level11_pos88_outg;
	wire node_level11_pos88_outp;
	neg_operator node_level11_pos88(.p1(p_in[88]), .g1(g_in[88]), .p0(node_level8_pos87_outp), .g0(node_level8_pos87_outg), .gp(node_level11_pos88_outg), .pp(node_level11_pos88_outp));
	wire node_level11_pos90_outg;
	wire node_level11_pos90_outp;
	neg_operator node_level11_pos90(.p1(p_in[90]), .g1(g_in[90]), .p0(node_level10_pos89_outp), .g0(node_level10_pos89_outg), .gp(node_level11_pos90_outg), .pp(node_level11_pos90_outp));
	wire node_level11_pos92_outg;
	wire node_level11_pos92_outp;
	neg_operator node_level11_pos92(.p1(p_in[92]), .g1(g_in[92]), .p0(~node_level9_pos91_outp), .g0(~node_level9_pos91_outg), .gp(node_level11_pos92_outg), .pp(node_level11_pos92_outp));
	wire node_level11_pos94_outg;
	wire node_level11_pos94_outp;
	neg_operator node_level11_pos94(.p1(p_in[94]), .g1(g_in[94]), .p0(node_level10_pos93_outp), .g0(node_level10_pos93_outg), .gp(node_level11_pos94_outg), .pp(node_level11_pos94_outp));
	wire node_level11_pos96_outg;
	wire node_level11_pos96_outp;
	neg_operator node_level11_pos96(.p1(p_in[96]), .g1(g_in[96]), .p0(~node_level7_pos95_outp), .g0(~node_level7_pos95_outg), .gp(node_level11_pos96_outg), .pp(node_level11_pos96_outp));
	wire node_level11_pos98_outg;
	wire node_level11_pos98_outp;
	neg_operator node_level11_pos98(.p1(p_in[98]), .g1(g_in[98]), .p0(node_level10_pos97_outp), .g0(node_level10_pos97_outg), .gp(node_level11_pos98_outg), .pp(node_level11_pos98_outp));
	wire node_level11_pos100_outg;
	wire node_level11_pos100_outp;
	neg_operator node_level11_pos100(.p1(p_in[100]), .g1(g_in[100]), .p0(~node_level9_pos99_outp), .g0(~node_level9_pos99_outg), .gp(node_level11_pos100_outg), .pp(node_level11_pos100_outp));
	wire node_level11_pos102_outg;
	wire node_level11_pos102_outp;
	neg_operator node_level11_pos102(.p1(p_in[102]), .g1(g_in[102]), .p0(node_level10_pos101_outp), .g0(node_level10_pos101_outg), .gp(node_level11_pos102_outg), .pp(node_level11_pos102_outp));
	wire node_level11_pos104_outg;
	wire node_level11_pos104_outp;
	neg_operator node_level11_pos104(.p1(p_in[104]), .g1(g_in[104]), .p0(node_level8_pos103_outp), .g0(node_level8_pos103_outg), .gp(node_level11_pos104_outg), .pp(node_level11_pos104_outp));
	wire node_level11_pos106_outg;
	wire node_level11_pos106_outp;
	neg_operator node_level11_pos106(.p1(p_in[106]), .g1(g_in[106]), .p0(node_level10_pos105_outp), .g0(node_level10_pos105_outg), .gp(node_level11_pos106_outg), .pp(node_level11_pos106_outp));
	wire node_level11_pos108_outg;
	wire node_level11_pos108_outp;
	neg_operator node_level11_pos108(.p1(p_in[108]), .g1(g_in[108]), .p0(~node_level9_pos107_outp), .g0(~node_level9_pos107_outg), .gp(node_level11_pos108_outg), .pp(node_level11_pos108_outp));
	wire node_level11_pos110_outg;
	wire node_level11_pos110_outp;
	neg_operator node_level11_pos110(.p1(p_in[110]), .g1(g_in[110]), .p0(node_level10_pos109_outp), .g0(node_level10_pos109_outg), .gp(node_level11_pos110_outg), .pp(node_level11_pos110_outp));
	wire node_level11_pos112_outg;
	wire node_level11_pos112_outp;
	neg_operator node_level11_pos112(.p1(p_in[112]), .g1(g_in[112]), .p0(~node_level7_pos111_outp), .g0(~node_level7_pos111_outg), .gp(node_level11_pos112_outg), .pp(node_level11_pos112_outp));
	wire node_level11_pos114_outg;
	wire node_level11_pos114_outp;
	neg_operator node_level11_pos114(.p1(p_in[114]), .g1(g_in[114]), .p0(node_level10_pos113_outp), .g0(node_level10_pos113_outg), .gp(node_level11_pos114_outg), .pp(node_level11_pos114_outp));
	wire node_level11_pos116_outg;
	wire node_level11_pos116_outp;
	neg_operator node_level11_pos116(.p1(p_in[116]), .g1(g_in[116]), .p0(~node_level9_pos115_outp), .g0(~node_level9_pos115_outg), .gp(node_level11_pos116_outg), .pp(node_level11_pos116_outp));
	wire node_level11_pos118_outg;
	wire node_level11_pos118_outp;
	neg_operator node_level11_pos118(.p1(p_in[118]), .g1(g_in[118]), .p0(node_level10_pos117_outp), .g0(node_level10_pos117_outg), .gp(node_level11_pos118_outg), .pp(node_level11_pos118_outp));
	wire node_level11_pos120_outg;
	wire node_level11_pos120_outp;
	neg_operator node_level11_pos120(.p1(p_in[120]), .g1(g_in[120]), .p0(node_level8_pos119_outp), .g0(node_level8_pos119_outg), .gp(node_level11_pos120_outg), .pp(node_level11_pos120_outp));
	wire node_level11_pos122_outg;
	wire node_level11_pos122_outp;
	neg_operator node_level11_pos122(.p1(p_in[122]), .g1(g_in[122]), .p0(node_level10_pos121_outp), .g0(node_level10_pos121_outg), .gp(node_level11_pos122_outg), .pp(node_level11_pos122_outp));
	wire node_level11_pos124_outg;
	wire node_level11_pos124_outp;
	neg_operator node_level11_pos124(.p1(p_in[124]), .g1(g_in[124]), .p0(~node_level9_pos123_outp), .g0(~node_level9_pos123_outg), .gp(node_level11_pos124_outg), .pp(node_level11_pos124_outp));
	wire node_level11_pos126_outg;
	wire node_level11_pos126_outp;
	neg_operator node_level11_pos126(.p1(p_in[126]), .g1(g_in[126]), .p0(node_level10_pos125_outp), .g0(node_level10_pos125_outg), .gp(node_level11_pos126_outg), .pp(node_level11_pos126_outp));


	assign s[0] = p_in[0];
	assign s[1] = p_in[1] ^ g_in[0];
	assign s[2] = p_in[2] ^ ~node_level1_pos1_outg;
	assign s[3] = p_in[3] ^ ~node_level11_pos2_outg;
	assign s[4] = p_in[4] ^ node_level2_pos3_outg;
	assign s[5] = p_in[5] ^ ~node_level11_pos4_outg;
	assign s[6] = p_in[6] ^ node_level10_pos5_outg;
	assign s[7] = p_in[7] ^ ~node_level11_pos6_outg;
	assign s[8] = p_in[8] ^ ~node_level3_pos7_outg;
	assign s[9] = p_in[9] ^ ~node_level11_pos8_outg;
	assign s[10] = p_in[10] ^ node_level10_pos9_outg;
	assign s[11] = p_in[11] ^ ~node_level11_pos10_outg;
	assign s[12] = p_in[12] ^ ~node_level9_pos11_outg;
	assign s[13] = p_in[13] ^ ~node_level11_pos12_outg;
	assign s[14] = p_in[14] ^ node_level10_pos13_outg;
	assign s[15] = p_in[15] ^ ~node_level11_pos14_outg;
	assign s[16] = p_in[16] ^ node_level4_pos15_outg;
	assign s[17] = p_in[17] ^ ~node_level11_pos16_outg;
	assign s[18] = p_in[18] ^ node_level10_pos17_outg;
	assign s[19] = p_in[19] ^ ~node_level11_pos18_outg;
	assign s[20] = p_in[20] ^ ~node_level9_pos19_outg;
	assign s[21] = p_in[21] ^ ~node_level11_pos20_outg;
	assign s[22] = p_in[22] ^ node_level10_pos21_outg;
	assign s[23] = p_in[23] ^ ~node_level11_pos22_outg;
	assign s[24] = p_in[24] ^ node_level8_pos23_outg;
	assign s[25] = p_in[25] ^ ~node_level11_pos24_outg;
	assign s[26] = p_in[26] ^ node_level10_pos25_outg;
	assign s[27] = p_in[27] ^ ~node_level11_pos26_outg;
	assign s[28] = p_in[28] ^ ~node_level9_pos27_outg;
	assign s[29] = p_in[29] ^ ~node_level11_pos28_outg;
	assign s[30] = p_in[30] ^ node_level10_pos29_outg;
	assign s[31] = p_in[31] ^ ~node_level11_pos30_outg;
	assign s[32] = p_in[32] ^ ~node_level5_pos31_outg;
	assign s[33] = p_in[33] ^ ~node_level11_pos32_outg;
	assign s[34] = p_in[34] ^ node_level10_pos33_outg;
	assign s[35] = p_in[35] ^ ~node_level11_pos34_outg;
	assign s[36] = p_in[36] ^ ~node_level9_pos35_outg;
	assign s[37] = p_in[37] ^ ~node_level11_pos36_outg;
	assign s[38] = p_in[38] ^ node_level10_pos37_outg;
	assign s[39] = p_in[39] ^ ~node_level11_pos38_outg;
	assign s[40] = p_in[40] ^ node_level8_pos39_outg;
	assign s[41] = p_in[41] ^ ~node_level11_pos40_outg;
	assign s[42] = p_in[42] ^ node_level10_pos41_outg;
	assign s[43] = p_in[43] ^ ~node_level11_pos42_outg;
	assign s[44] = p_in[44] ^ ~node_level9_pos43_outg;
	assign s[45] = p_in[45] ^ ~node_level11_pos44_outg;
	assign s[46] = p_in[46] ^ node_level10_pos45_outg;
	assign s[47] = p_in[47] ^ ~node_level11_pos46_outg;
	assign s[48] = p_in[48] ^ node_level6_pos47_outg;
	assign s[49] = p_in[49] ^ ~node_level11_pos48_outg;
	assign s[50] = p_in[50] ^ node_level10_pos49_outg;
	assign s[51] = p_in[51] ^ ~node_level11_pos50_outg;
	assign s[52] = p_in[52] ^ ~node_level9_pos51_outg;
	assign s[53] = p_in[53] ^ ~node_level11_pos52_outg;
	assign s[54] = p_in[54] ^ node_level10_pos53_outg;
	assign s[55] = p_in[55] ^ ~node_level11_pos54_outg;
	assign s[56] = p_in[56] ^ node_level8_pos55_outg;
	assign s[57] = p_in[57] ^ ~node_level11_pos56_outg;
	assign s[58] = p_in[58] ^ node_level10_pos57_outg;
	assign s[59] = p_in[59] ^ ~node_level11_pos58_outg;
	assign s[60] = p_in[60] ^ ~node_level9_pos59_outg;
	assign s[61] = p_in[61] ^ ~node_level11_pos60_outg;
	assign s[62] = p_in[62] ^ node_level10_pos61_outg;
	assign s[63] = p_in[63] ^ ~node_level11_pos62_outg;
	assign s[64] = p_in[64] ^ node_level6_pos63_outg;
	assign s[65] = p_in[65] ^ ~node_level11_pos64_outg;
	assign s[66] = p_in[66] ^ node_level10_pos65_outg;
	assign s[67] = p_in[67] ^ ~node_level11_pos66_outg;
	assign s[68] = p_in[68] ^ ~node_level9_pos67_outg;
	assign s[69] = p_in[69] ^ ~node_level11_pos68_outg;
	assign s[70] = p_in[70] ^ node_level10_pos69_outg;
	assign s[71] = p_in[71] ^ ~node_level11_pos70_outg;
	assign s[72] = p_in[72] ^ node_level8_pos71_outg;
	assign s[73] = p_in[73] ^ ~node_level11_pos72_outg;
	assign s[74] = p_in[74] ^ node_level10_pos73_outg;
	assign s[75] = p_in[75] ^ ~node_level11_pos74_outg;
	assign s[76] = p_in[76] ^ ~node_level9_pos75_outg;
	assign s[77] = p_in[77] ^ ~node_level11_pos76_outg;
	assign s[78] = p_in[78] ^ node_level10_pos77_outg;
	assign s[79] = p_in[79] ^ ~node_level11_pos78_outg;
	assign s[80] = p_in[80] ^ ~node_level7_pos79_outg;
	assign s[81] = p_in[81] ^ ~node_level11_pos80_outg;
	assign s[82] = p_in[82] ^ node_level10_pos81_outg;
	assign s[83] = p_in[83] ^ ~node_level11_pos82_outg;
	assign s[84] = p_in[84] ^ ~node_level9_pos83_outg;
	assign s[85] = p_in[85] ^ ~node_level11_pos84_outg;
	assign s[86] = p_in[86] ^ node_level10_pos85_outg;
	assign s[87] = p_in[87] ^ ~node_level11_pos86_outg;
	assign s[88] = p_in[88] ^ node_level8_pos87_outg;
	assign s[89] = p_in[89] ^ ~node_level11_pos88_outg;
	assign s[90] = p_in[90] ^ node_level10_pos89_outg;
	assign s[91] = p_in[91] ^ ~node_level11_pos90_outg;
	assign s[92] = p_in[92] ^ ~node_level9_pos91_outg;
	assign s[93] = p_in[93] ^ ~node_level11_pos92_outg;
	assign s[94] = p_in[94] ^ node_level10_pos93_outg;
	assign s[95] = p_in[95] ^ ~node_level11_pos94_outg;
	assign s[96] = p_in[96] ^ ~node_level7_pos95_outg;
	assign s[97] = p_in[97] ^ ~node_level11_pos96_outg;
	assign s[98] = p_in[98] ^ node_level10_pos97_outg;
	assign s[99] = p_in[99] ^ ~node_level11_pos98_outg;
	assign s[100] = p_in[100] ^ ~node_level9_pos99_outg;
	assign s[101] = p_in[101] ^ ~node_level11_pos100_outg;
	assign s[102] = p_in[102] ^ node_level10_pos101_outg;
	assign s[103] = p_in[103] ^ ~node_level11_pos102_outg;
	assign s[104] = p_in[104] ^ node_level8_pos103_outg;
	assign s[105] = p_in[105] ^ ~node_level11_pos104_outg;
	assign s[106] = p_in[106] ^ node_level10_pos105_outg;
	assign s[107] = p_in[107] ^ ~node_level11_pos106_outg;
	assign s[108] = p_in[108] ^ ~node_level9_pos107_outg;
	assign s[109] = p_in[109] ^ ~node_level11_pos108_outg;
	assign s[110] = p_in[110] ^ node_level10_pos109_outg;
	assign s[111] = p_in[111] ^ ~node_level11_pos110_outg;
	assign s[112] = p_in[112] ^ ~node_level7_pos111_outg;
	assign s[113] = p_in[113] ^ ~node_level11_pos112_outg;
	assign s[114] = p_in[114] ^ node_level10_pos113_outg;
	assign s[115] = p_in[115] ^ ~node_level11_pos114_outg;
	assign s[116] = p_in[116] ^ ~node_level9_pos115_outg;
	assign s[117] = p_in[117] ^ ~node_level11_pos116_outg;
	assign s[118] = p_in[118] ^ node_level10_pos117_outg;
	assign s[119] = p_in[119] ^ ~node_level11_pos118_outg;
	assign s[120] = p_in[120] ^ node_level8_pos119_outg;
	assign s[121] = p_in[121] ^ ~node_level11_pos120_outg;
	assign s[122] = p_in[122] ^ node_level10_pos121_outg;
	assign s[123] = p_in[123] ^ ~node_level11_pos122_outg;
	assign s[124] = p_in[124] ^ ~node_level9_pos123_outg;
	assign s[125] = p_in[125] ^ ~node_level11_pos124_outg;
	assign s[126] = p_in[126] ^ node_level10_pos125_outg;
	assign s[127] = p_in[127] ^ ~node_level11_pos126_outg;
	// AND count: 169, NAND count: 253, OR count: 84, NOR count: 253, NOT count: 84, Transistor count: 4724
endmodule

