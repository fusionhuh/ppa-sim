`ifndef CARRY_OPERATOR
`include "carry_operator.v"
`endif
`ifndef NEG_CARRY_OPERATOR
`include "neg_operator.v"
`endif
`ifndef POS_CARRY_OPERATOR
`include "pos_operator.v"
`endif
`define KS32
// number of levels: 6
// number of nodes: 129
// NAND count: 129, AND count: 75
// NOR count: 129, OR count: 54
// NOT count: 41, Transistor count: 1888
module ks32(x1, x2, s, cin, cout, p_out, g_out);
	input[31:0]x1;
	input[31:0]x2;
	input cin;
	wire[31:0]p_in;
	wire[31:0]g_in;
	output[31:0]s;
	output cout;

	output[31:0]p_out;
	output[31:0]g_out;
	assign p_in = x1 ^ x2;
	assign p_out = p_in;
	assign g_in[31:1] = x1[31:1] & x2[31:1];
	assign g_in[0] = (x1[0] & x2[0]) | (p_in[0] & cin);
	assign g_out = g_in;
	wire node_level1_pos1_outg;
	wire node_level1_pos1_outp;
	neg_operator node_level1_pos1(.p1(p_in[1]), .g1(g_in[1]), .p0(p_in[0]), .g0(g_in[0]), .gp(node_level1_pos1_outg), .pp(node_level1_pos1_outp));
	wire node_level1_pos2_outg;
	wire node_level1_pos2_outp;
	neg_operator node_level1_pos2(.p1(p_in[2]), .g1(g_in[2]), .p0(p_in[1]), .g0(g_in[1]), .gp(node_level1_pos2_outg), .pp(node_level1_pos2_outp));
	wire node_level1_pos3_outg;
	wire node_level1_pos3_outp;
	neg_operator node_level1_pos3(.p1(p_in[3]), .g1(g_in[3]), .p0(p_in[2]), .g0(g_in[2]), .gp(node_level1_pos3_outg), .pp(node_level1_pos3_outp));
	wire node_level1_pos4_outg;
	wire node_level1_pos4_outp;
	neg_operator node_level1_pos4(.p1(p_in[4]), .g1(g_in[4]), .p0(p_in[3]), .g0(g_in[3]), .gp(node_level1_pos4_outg), .pp(node_level1_pos4_outp));
	wire node_level1_pos5_outg;
	wire node_level1_pos5_outp;
	neg_operator node_level1_pos5(.p1(p_in[5]), .g1(g_in[5]), .p0(p_in[4]), .g0(g_in[4]), .gp(node_level1_pos5_outg), .pp(node_level1_pos5_outp));
	wire node_level1_pos6_outg;
	wire node_level1_pos6_outp;
	neg_operator node_level1_pos6(.p1(p_in[6]), .g1(g_in[6]), .p0(p_in[5]), .g0(g_in[5]), .gp(node_level1_pos6_outg), .pp(node_level1_pos6_outp));
	wire node_level1_pos7_outg;
	wire node_level1_pos7_outp;
	neg_operator node_level1_pos7(.p1(p_in[7]), .g1(g_in[7]), .p0(p_in[6]), .g0(g_in[6]), .gp(node_level1_pos7_outg), .pp(node_level1_pos7_outp));
	wire node_level1_pos8_outg;
	wire node_level1_pos8_outp;
	neg_operator node_level1_pos8(.p1(p_in[8]), .g1(g_in[8]), .p0(p_in[7]), .g0(g_in[7]), .gp(node_level1_pos8_outg), .pp(node_level1_pos8_outp));
	wire node_level1_pos9_outg;
	wire node_level1_pos9_outp;
	neg_operator node_level1_pos9(.p1(p_in[9]), .g1(g_in[9]), .p0(p_in[8]), .g0(g_in[8]), .gp(node_level1_pos9_outg), .pp(node_level1_pos9_outp));
	wire node_level1_pos10_outg;
	wire node_level1_pos10_outp;
	neg_operator node_level1_pos10(.p1(p_in[10]), .g1(g_in[10]), .p0(p_in[9]), .g0(g_in[9]), .gp(node_level1_pos10_outg), .pp(node_level1_pos10_outp));
	wire node_level1_pos11_outg;
	wire node_level1_pos11_outp;
	neg_operator node_level1_pos11(.p1(p_in[11]), .g1(g_in[11]), .p0(p_in[10]), .g0(g_in[10]), .gp(node_level1_pos11_outg), .pp(node_level1_pos11_outp));
	wire node_level1_pos12_outg;
	wire node_level1_pos12_outp;
	neg_operator node_level1_pos12(.p1(p_in[12]), .g1(g_in[12]), .p0(p_in[11]), .g0(g_in[11]), .gp(node_level1_pos12_outg), .pp(node_level1_pos12_outp));
	wire node_level1_pos13_outg;
	wire node_level1_pos13_outp;
	neg_operator node_level1_pos13(.p1(p_in[13]), .g1(g_in[13]), .p0(p_in[12]), .g0(g_in[12]), .gp(node_level1_pos13_outg), .pp(node_level1_pos13_outp));
	wire node_level1_pos14_outg;
	wire node_level1_pos14_outp;
	neg_operator node_level1_pos14(.p1(p_in[14]), .g1(g_in[14]), .p0(p_in[13]), .g0(g_in[13]), .gp(node_level1_pos14_outg), .pp(node_level1_pos14_outp));
	wire node_level1_pos15_outg;
	wire node_level1_pos15_outp;
	neg_operator node_level1_pos15(.p1(p_in[15]), .g1(g_in[15]), .p0(p_in[14]), .g0(g_in[14]), .gp(node_level1_pos15_outg), .pp(node_level1_pos15_outp));
	wire node_level1_pos16_outg;
	wire node_level1_pos16_outp;
	neg_operator node_level1_pos16(.p1(p_in[16]), .g1(g_in[16]), .p0(p_in[15]), .g0(g_in[15]), .gp(node_level1_pos16_outg), .pp(node_level1_pos16_outp));
	wire node_level1_pos17_outg;
	wire node_level1_pos17_outp;
	neg_operator node_level1_pos17(.p1(p_in[17]), .g1(g_in[17]), .p0(p_in[16]), .g0(g_in[16]), .gp(node_level1_pos17_outg), .pp(node_level1_pos17_outp));
	wire node_level1_pos18_outg;
	wire node_level1_pos18_outp;
	neg_operator node_level1_pos18(.p1(p_in[18]), .g1(g_in[18]), .p0(p_in[17]), .g0(g_in[17]), .gp(node_level1_pos18_outg), .pp(node_level1_pos18_outp));
	wire node_level1_pos19_outg;
	wire node_level1_pos19_outp;
	neg_operator node_level1_pos19(.p1(p_in[19]), .g1(g_in[19]), .p0(p_in[18]), .g0(g_in[18]), .gp(node_level1_pos19_outg), .pp(node_level1_pos19_outp));
	wire node_level1_pos20_outg;
	wire node_level1_pos20_outp;
	neg_operator node_level1_pos20(.p1(p_in[20]), .g1(g_in[20]), .p0(p_in[19]), .g0(g_in[19]), .gp(node_level1_pos20_outg), .pp(node_level1_pos20_outp));
	wire node_level1_pos21_outg;
	wire node_level1_pos21_outp;
	neg_operator node_level1_pos21(.p1(p_in[21]), .g1(g_in[21]), .p0(p_in[20]), .g0(g_in[20]), .gp(node_level1_pos21_outg), .pp(node_level1_pos21_outp));
	wire node_level1_pos22_outg;
	wire node_level1_pos22_outp;
	neg_operator node_level1_pos22(.p1(p_in[22]), .g1(g_in[22]), .p0(p_in[21]), .g0(g_in[21]), .gp(node_level1_pos22_outg), .pp(node_level1_pos22_outp));
	wire node_level1_pos23_outg;
	wire node_level1_pos23_outp;
	neg_operator node_level1_pos23(.p1(p_in[23]), .g1(g_in[23]), .p0(p_in[22]), .g0(g_in[22]), .gp(node_level1_pos23_outg), .pp(node_level1_pos23_outp));
	wire node_level1_pos24_outg;
	wire node_level1_pos24_outp;
	neg_operator node_level1_pos24(.p1(p_in[24]), .g1(g_in[24]), .p0(p_in[23]), .g0(g_in[23]), .gp(node_level1_pos24_outg), .pp(node_level1_pos24_outp));
	wire node_level1_pos25_outg;
	wire node_level1_pos25_outp;
	neg_operator node_level1_pos25(.p1(p_in[25]), .g1(g_in[25]), .p0(p_in[24]), .g0(g_in[24]), .gp(node_level1_pos25_outg), .pp(node_level1_pos25_outp));
	wire node_level1_pos26_outg;
	wire node_level1_pos26_outp;
	neg_operator node_level1_pos26(.p1(p_in[26]), .g1(g_in[26]), .p0(p_in[25]), .g0(g_in[25]), .gp(node_level1_pos26_outg), .pp(node_level1_pos26_outp));
	wire node_level1_pos27_outg;
	wire node_level1_pos27_outp;
	neg_operator node_level1_pos27(.p1(p_in[27]), .g1(g_in[27]), .p0(p_in[26]), .g0(g_in[26]), .gp(node_level1_pos27_outg), .pp(node_level1_pos27_outp));
	wire node_level1_pos28_outg;
	wire node_level1_pos28_outp;
	neg_operator node_level1_pos28(.p1(p_in[28]), .g1(g_in[28]), .p0(p_in[27]), .g0(g_in[27]), .gp(node_level1_pos28_outg), .pp(node_level1_pos28_outp));
	wire node_level1_pos29_outg;
	wire node_level1_pos29_outp;
	neg_operator node_level1_pos29(.p1(p_in[29]), .g1(g_in[29]), .p0(p_in[28]), .g0(g_in[28]), .gp(node_level1_pos29_outg), .pp(node_level1_pos29_outp));
	wire node_level1_pos30_outg;
	wire node_level1_pos30_outp;
	neg_operator node_level1_pos30(.p1(p_in[30]), .g1(g_in[30]), .p0(p_in[29]), .g0(g_in[29]), .gp(node_level1_pos30_outg), .pp(node_level1_pos30_outp));
	wire node_level1_pos31_outg;
	wire node_level1_pos31_outp;
	neg_operator node_level1_pos31(.p1(p_in[31]), .g1(g_in[31]), .p0(p_in[30]), .g0(g_in[30]), .gp(node_level1_pos31_outg), .pp(node_level1_pos31_outp));
	wire node_level2_pos2_outg;
	wire node_level2_pos2_outp;
	pos_operator node_level2_pos2(.p1(node_level1_pos2_outp), .g1(node_level1_pos2_outg), .p0(~p_in[0]), .g0(~g_in[0]), .gp(node_level2_pos2_outg), .pp(node_level2_pos2_outp));
	wire node_level2_pos3_outg;
	wire node_level2_pos3_outp;
	pos_operator node_level2_pos3(.p1(node_level1_pos3_outp), .g1(node_level1_pos3_outg), .p0(node_level1_pos1_outp), .g0(node_level1_pos1_outg), .gp(node_level2_pos3_outg), .pp(node_level2_pos3_outp));
	wire node_level2_pos4_outg;
	wire node_level2_pos4_outp;
	pos_operator node_level2_pos4(.p1(node_level1_pos4_outp), .g1(node_level1_pos4_outg), .p0(node_level1_pos2_outp), .g0(node_level1_pos2_outg), .gp(node_level2_pos4_outg), .pp(node_level2_pos4_outp));
	wire node_level2_pos5_outg;
	wire node_level2_pos5_outp;
	pos_operator node_level2_pos5(.p1(node_level1_pos5_outp), .g1(node_level1_pos5_outg), .p0(node_level1_pos3_outp), .g0(node_level1_pos3_outg), .gp(node_level2_pos5_outg), .pp(node_level2_pos5_outp));
	wire node_level2_pos6_outg;
	wire node_level2_pos6_outp;
	pos_operator node_level2_pos6(.p1(node_level1_pos6_outp), .g1(node_level1_pos6_outg), .p0(node_level1_pos4_outp), .g0(node_level1_pos4_outg), .gp(node_level2_pos6_outg), .pp(node_level2_pos6_outp));
	wire node_level2_pos7_outg;
	wire node_level2_pos7_outp;
	pos_operator node_level2_pos7(.p1(node_level1_pos7_outp), .g1(node_level1_pos7_outg), .p0(node_level1_pos5_outp), .g0(node_level1_pos5_outg), .gp(node_level2_pos7_outg), .pp(node_level2_pos7_outp));
	wire node_level2_pos8_outg;
	wire node_level2_pos8_outp;
	pos_operator node_level2_pos8(.p1(node_level1_pos8_outp), .g1(node_level1_pos8_outg), .p0(node_level1_pos6_outp), .g0(node_level1_pos6_outg), .gp(node_level2_pos8_outg), .pp(node_level2_pos8_outp));
	wire node_level2_pos9_outg;
	wire node_level2_pos9_outp;
	pos_operator node_level2_pos9(.p1(node_level1_pos9_outp), .g1(node_level1_pos9_outg), .p0(node_level1_pos7_outp), .g0(node_level1_pos7_outg), .gp(node_level2_pos9_outg), .pp(node_level2_pos9_outp));
	wire node_level2_pos10_outg;
	wire node_level2_pos10_outp;
	pos_operator node_level2_pos10(.p1(node_level1_pos10_outp), .g1(node_level1_pos10_outg), .p0(node_level1_pos8_outp), .g0(node_level1_pos8_outg), .gp(node_level2_pos10_outg), .pp(node_level2_pos10_outp));
	wire node_level2_pos11_outg;
	wire node_level2_pos11_outp;
	pos_operator node_level2_pos11(.p1(node_level1_pos11_outp), .g1(node_level1_pos11_outg), .p0(node_level1_pos9_outp), .g0(node_level1_pos9_outg), .gp(node_level2_pos11_outg), .pp(node_level2_pos11_outp));
	wire node_level2_pos12_outg;
	wire node_level2_pos12_outp;
	pos_operator node_level2_pos12(.p1(node_level1_pos12_outp), .g1(node_level1_pos12_outg), .p0(node_level1_pos10_outp), .g0(node_level1_pos10_outg), .gp(node_level2_pos12_outg), .pp(node_level2_pos12_outp));
	wire node_level2_pos13_outg;
	wire node_level2_pos13_outp;
	pos_operator node_level2_pos13(.p1(node_level1_pos13_outp), .g1(node_level1_pos13_outg), .p0(node_level1_pos11_outp), .g0(node_level1_pos11_outg), .gp(node_level2_pos13_outg), .pp(node_level2_pos13_outp));
	wire node_level2_pos14_outg;
	wire node_level2_pos14_outp;
	pos_operator node_level2_pos14(.p1(node_level1_pos14_outp), .g1(node_level1_pos14_outg), .p0(node_level1_pos12_outp), .g0(node_level1_pos12_outg), .gp(node_level2_pos14_outg), .pp(node_level2_pos14_outp));
	wire node_level2_pos15_outg;
	wire node_level2_pos15_outp;
	pos_operator node_level2_pos15(.p1(node_level1_pos15_outp), .g1(node_level1_pos15_outg), .p0(node_level1_pos13_outp), .g0(node_level1_pos13_outg), .gp(node_level2_pos15_outg), .pp(node_level2_pos15_outp));
	wire node_level2_pos16_outg;
	wire node_level2_pos16_outp;
	pos_operator node_level2_pos16(.p1(node_level1_pos16_outp), .g1(node_level1_pos16_outg), .p0(node_level1_pos14_outp), .g0(node_level1_pos14_outg), .gp(node_level2_pos16_outg), .pp(node_level2_pos16_outp));
	wire node_level2_pos17_outg;
	wire node_level2_pos17_outp;
	pos_operator node_level2_pos17(.p1(node_level1_pos17_outp), .g1(node_level1_pos17_outg), .p0(node_level1_pos15_outp), .g0(node_level1_pos15_outg), .gp(node_level2_pos17_outg), .pp(node_level2_pos17_outp));
	wire node_level2_pos18_outg;
	wire node_level2_pos18_outp;
	pos_operator node_level2_pos18(.p1(node_level1_pos18_outp), .g1(node_level1_pos18_outg), .p0(node_level1_pos16_outp), .g0(node_level1_pos16_outg), .gp(node_level2_pos18_outg), .pp(node_level2_pos18_outp));
	wire node_level2_pos19_outg;
	wire node_level2_pos19_outp;
	pos_operator node_level2_pos19(.p1(node_level1_pos19_outp), .g1(node_level1_pos19_outg), .p0(node_level1_pos17_outp), .g0(node_level1_pos17_outg), .gp(node_level2_pos19_outg), .pp(node_level2_pos19_outp));
	wire node_level2_pos20_outg;
	wire node_level2_pos20_outp;
	pos_operator node_level2_pos20(.p1(node_level1_pos20_outp), .g1(node_level1_pos20_outg), .p0(node_level1_pos18_outp), .g0(node_level1_pos18_outg), .gp(node_level2_pos20_outg), .pp(node_level2_pos20_outp));
	wire node_level2_pos21_outg;
	wire node_level2_pos21_outp;
	pos_operator node_level2_pos21(.p1(node_level1_pos21_outp), .g1(node_level1_pos21_outg), .p0(node_level1_pos19_outp), .g0(node_level1_pos19_outg), .gp(node_level2_pos21_outg), .pp(node_level2_pos21_outp));
	wire node_level2_pos22_outg;
	wire node_level2_pos22_outp;
	pos_operator node_level2_pos22(.p1(node_level1_pos22_outp), .g1(node_level1_pos22_outg), .p0(node_level1_pos20_outp), .g0(node_level1_pos20_outg), .gp(node_level2_pos22_outg), .pp(node_level2_pos22_outp));
	wire node_level2_pos23_outg;
	wire node_level2_pos23_outp;
	pos_operator node_level2_pos23(.p1(node_level1_pos23_outp), .g1(node_level1_pos23_outg), .p0(node_level1_pos21_outp), .g0(node_level1_pos21_outg), .gp(node_level2_pos23_outg), .pp(node_level2_pos23_outp));
	wire node_level2_pos24_outg;
	wire node_level2_pos24_outp;
	pos_operator node_level2_pos24(.p1(node_level1_pos24_outp), .g1(node_level1_pos24_outg), .p0(node_level1_pos22_outp), .g0(node_level1_pos22_outg), .gp(node_level2_pos24_outg), .pp(node_level2_pos24_outp));
	wire node_level2_pos25_outg;
	wire node_level2_pos25_outp;
	pos_operator node_level2_pos25(.p1(node_level1_pos25_outp), .g1(node_level1_pos25_outg), .p0(node_level1_pos23_outp), .g0(node_level1_pos23_outg), .gp(node_level2_pos25_outg), .pp(node_level2_pos25_outp));
	wire node_level2_pos26_outg;
	wire node_level2_pos26_outp;
	pos_operator node_level2_pos26(.p1(node_level1_pos26_outp), .g1(node_level1_pos26_outg), .p0(node_level1_pos24_outp), .g0(node_level1_pos24_outg), .gp(node_level2_pos26_outg), .pp(node_level2_pos26_outp));
	wire node_level2_pos27_outg;
	wire node_level2_pos27_outp;
	pos_operator node_level2_pos27(.p1(node_level1_pos27_outp), .g1(node_level1_pos27_outg), .p0(node_level1_pos25_outp), .g0(node_level1_pos25_outg), .gp(node_level2_pos27_outg), .pp(node_level2_pos27_outp));
	wire node_level2_pos28_outg;
	wire node_level2_pos28_outp;
	pos_operator node_level2_pos28(.p1(node_level1_pos28_outp), .g1(node_level1_pos28_outg), .p0(node_level1_pos26_outp), .g0(node_level1_pos26_outg), .gp(node_level2_pos28_outg), .pp(node_level2_pos28_outp));
	wire node_level2_pos29_outg;
	wire node_level2_pos29_outp;
	pos_operator node_level2_pos29(.p1(node_level1_pos29_outp), .g1(node_level1_pos29_outg), .p0(node_level1_pos27_outp), .g0(node_level1_pos27_outg), .gp(node_level2_pos29_outg), .pp(node_level2_pos29_outp));
	wire node_level2_pos30_outg;
	wire node_level2_pos30_outp;
	pos_operator node_level2_pos30(.p1(node_level1_pos30_outp), .g1(node_level1_pos30_outg), .p0(node_level1_pos28_outp), .g0(node_level1_pos28_outg), .gp(node_level2_pos30_outg), .pp(node_level2_pos30_outp));
	wire node_level2_pos31_outg;
	wire node_level2_pos31_outp;
	pos_operator node_level2_pos31(.p1(node_level1_pos31_outp), .g1(node_level1_pos31_outg), .p0(node_level1_pos29_outp), .g0(node_level1_pos29_outg), .gp(node_level2_pos31_outg), .pp(node_level2_pos31_outp));
	wire node_level3_pos4_outg;
	wire node_level3_pos4_outp;
	neg_operator node_level3_pos4(.p1(node_level2_pos4_outp), .g1(node_level2_pos4_outg), .p0(p_in[0]), .g0(g_in[0]), .gp(node_level3_pos4_outg), .pp(node_level3_pos4_outp));
	wire node_level3_pos5_outg;
	wire node_level3_pos5_outp;
	neg_operator node_level3_pos5(.p1(node_level2_pos5_outp), .g1(node_level2_pos5_outg), .p0(~node_level1_pos1_outp), .g0(~node_level1_pos1_outg), .gp(node_level3_pos5_outg), .pp(node_level3_pos5_outp));
	wire node_level3_pos6_outg;
	wire node_level3_pos6_outp;
	neg_operator node_level3_pos6(.p1(node_level2_pos6_outp), .g1(node_level2_pos6_outg), .p0(node_level2_pos2_outp), .g0(node_level2_pos2_outg), .gp(node_level3_pos6_outg), .pp(node_level3_pos6_outp));
	wire node_level3_pos7_outg;
	wire node_level3_pos7_outp;
	neg_operator node_level3_pos7(.p1(node_level2_pos7_outp), .g1(node_level2_pos7_outg), .p0(node_level2_pos3_outp), .g0(node_level2_pos3_outg), .gp(node_level3_pos7_outg), .pp(node_level3_pos7_outp));
	wire node_level3_pos8_outg;
	wire node_level3_pos8_outp;
	neg_operator node_level3_pos8(.p1(node_level2_pos8_outp), .g1(node_level2_pos8_outg), .p0(node_level2_pos4_outp), .g0(node_level2_pos4_outg), .gp(node_level3_pos8_outg), .pp(node_level3_pos8_outp));
	wire node_level3_pos9_outg;
	wire node_level3_pos9_outp;
	neg_operator node_level3_pos9(.p1(node_level2_pos9_outp), .g1(node_level2_pos9_outg), .p0(node_level2_pos5_outp), .g0(node_level2_pos5_outg), .gp(node_level3_pos9_outg), .pp(node_level3_pos9_outp));
	wire node_level3_pos10_outg;
	wire node_level3_pos10_outp;
	neg_operator node_level3_pos10(.p1(node_level2_pos10_outp), .g1(node_level2_pos10_outg), .p0(node_level2_pos6_outp), .g0(node_level2_pos6_outg), .gp(node_level3_pos10_outg), .pp(node_level3_pos10_outp));
	wire node_level3_pos11_outg;
	wire node_level3_pos11_outp;
	neg_operator node_level3_pos11(.p1(node_level2_pos11_outp), .g1(node_level2_pos11_outg), .p0(node_level2_pos7_outp), .g0(node_level2_pos7_outg), .gp(node_level3_pos11_outg), .pp(node_level3_pos11_outp));
	wire node_level3_pos12_outg;
	wire node_level3_pos12_outp;
	neg_operator node_level3_pos12(.p1(node_level2_pos12_outp), .g1(node_level2_pos12_outg), .p0(node_level2_pos8_outp), .g0(node_level2_pos8_outg), .gp(node_level3_pos12_outg), .pp(node_level3_pos12_outp));
	wire node_level3_pos13_outg;
	wire node_level3_pos13_outp;
	neg_operator node_level3_pos13(.p1(node_level2_pos13_outp), .g1(node_level2_pos13_outg), .p0(node_level2_pos9_outp), .g0(node_level2_pos9_outg), .gp(node_level3_pos13_outg), .pp(node_level3_pos13_outp));
	wire node_level3_pos14_outg;
	wire node_level3_pos14_outp;
	neg_operator node_level3_pos14(.p1(node_level2_pos14_outp), .g1(node_level2_pos14_outg), .p0(node_level2_pos10_outp), .g0(node_level2_pos10_outg), .gp(node_level3_pos14_outg), .pp(node_level3_pos14_outp));
	wire node_level3_pos15_outg;
	wire node_level3_pos15_outp;
	neg_operator node_level3_pos15(.p1(node_level2_pos15_outp), .g1(node_level2_pos15_outg), .p0(node_level2_pos11_outp), .g0(node_level2_pos11_outg), .gp(node_level3_pos15_outg), .pp(node_level3_pos15_outp));
	wire node_level3_pos16_outg;
	wire node_level3_pos16_outp;
	neg_operator node_level3_pos16(.p1(node_level2_pos16_outp), .g1(node_level2_pos16_outg), .p0(node_level2_pos12_outp), .g0(node_level2_pos12_outg), .gp(node_level3_pos16_outg), .pp(node_level3_pos16_outp));
	wire node_level3_pos17_outg;
	wire node_level3_pos17_outp;
	neg_operator node_level3_pos17(.p1(node_level2_pos17_outp), .g1(node_level2_pos17_outg), .p0(node_level2_pos13_outp), .g0(node_level2_pos13_outg), .gp(node_level3_pos17_outg), .pp(node_level3_pos17_outp));
	wire node_level3_pos18_outg;
	wire node_level3_pos18_outp;
	neg_operator node_level3_pos18(.p1(node_level2_pos18_outp), .g1(node_level2_pos18_outg), .p0(node_level2_pos14_outp), .g0(node_level2_pos14_outg), .gp(node_level3_pos18_outg), .pp(node_level3_pos18_outp));
	wire node_level3_pos19_outg;
	wire node_level3_pos19_outp;
	neg_operator node_level3_pos19(.p1(node_level2_pos19_outp), .g1(node_level2_pos19_outg), .p0(node_level2_pos15_outp), .g0(node_level2_pos15_outg), .gp(node_level3_pos19_outg), .pp(node_level3_pos19_outp));
	wire node_level3_pos20_outg;
	wire node_level3_pos20_outp;
	neg_operator node_level3_pos20(.p1(node_level2_pos20_outp), .g1(node_level2_pos20_outg), .p0(node_level2_pos16_outp), .g0(node_level2_pos16_outg), .gp(node_level3_pos20_outg), .pp(node_level3_pos20_outp));
	wire node_level3_pos21_outg;
	wire node_level3_pos21_outp;
	neg_operator node_level3_pos21(.p1(node_level2_pos21_outp), .g1(node_level2_pos21_outg), .p0(node_level2_pos17_outp), .g0(node_level2_pos17_outg), .gp(node_level3_pos21_outg), .pp(node_level3_pos21_outp));
	wire node_level3_pos22_outg;
	wire node_level3_pos22_outp;
	neg_operator node_level3_pos22(.p1(node_level2_pos22_outp), .g1(node_level2_pos22_outg), .p0(node_level2_pos18_outp), .g0(node_level2_pos18_outg), .gp(node_level3_pos22_outg), .pp(node_level3_pos22_outp));
	wire node_level3_pos23_outg;
	wire node_level3_pos23_outp;
	neg_operator node_level3_pos23(.p1(node_level2_pos23_outp), .g1(node_level2_pos23_outg), .p0(node_level2_pos19_outp), .g0(node_level2_pos19_outg), .gp(node_level3_pos23_outg), .pp(node_level3_pos23_outp));
	wire node_level3_pos24_outg;
	wire node_level3_pos24_outp;
	neg_operator node_level3_pos24(.p1(node_level2_pos24_outp), .g1(node_level2_pos24_outg), .p0(node_level2_pos20_outp), .g0(node_level2_pos20_outg), .gp(node_level3_pos24_outg), .pp(node_level3_pos24_outp));
	wire node_level3_pos25_outg;
	wire node_level3_pos25_outp;
	neg_operator node_level3_pos25(.p1(node_level2_pos25_outp), .g1(node_level2_pos25_outg), .p0(node_level2_pos21_outp), .g0(node_level2_pos21_outg), .gp(node_level3_pos25_outg), .pp(node_level3_pos25_outp));
	wire node_level3_pos26_outg;
	wire node_level3_pos26_outp;
	neg_operator node_level3_pos26(.p1(node_level2_pos26_outp), .g1(node_level2_pos26_outg), .p0(node_level2_pos22_outp), .g0(node_level2_pos22_outg), .gp(node_level3_pos26_outg), .pp(node_level3_pos26_outp));
	wire node_level3_pos27_outg;
	wire node_level3_pos27_outp;
	neg_operator node_level3_pos27(.p1(node_level2_pos27_outp), .g1(node_level2_pos27_outg), .p0(node_level2_pos23_outp), .g0(node_level2_pos23_outg), .gp(node_level3_pos27_outg), .pp(node_level3_pos27_outp));
	wire node_level3_pos28_outg;
	wire node_level3_pos28_outp;
	neg_operator node_level3_pos28(.p1(node_level2_pos28_outp), .g1(node_level2_pos28_outg), .p0(node_level2_pos24_outp), .g0(node_level2_pos24_outg), .gp(node_level3_pos28_outg), .pp(node_level3_pos28_outp));
	wire node_level3_pos29_outg;
	wire node_level3_pos29_outp;
	neg_operator node_level3_pos29(.p1(node_level2_pos29_outp), .g1(node_level2_pos29_outg), .p0(node_level2_pos25_outp), .g0(node_level2_pos25_outg), .gp(node_level3_pos29_outg), .pp(node_level3_pos29_outp));
	wire node_level3_pos30_outg;
	wire node_level3_pos30_outp;
	neg_operator node_level3_pos30(.p1(node_level2_pos30_outp), .g1(node_level2_pos30_outg), .p0(node_level2_pos26_outp), .g0(node_level2_pos26_outg), .gp(node_level3_pos30_outg), .pp(node_level3_pos30_outp));
	wire node_level3_pos31_outg;
	wire node_level3_pos31_outp;
	neg_operator node_level3_pos31(.p1(node_level2_pos31_outp), .g1(node_level2_pos31_outg), .p0(node_level2_pos27_outp), .g0(node_level2_pos27_outg), .gp(node_level3_pos31_outg), .pp(node_level3_pos31_outp));
	wire node_level4_pos8_outg;
	wire node_level4_pos8_outp;
	pos_operator node_level4_pos8(.p1(node_level3_pos8_outp), .g1(node_level3_pos8_outg), .p0(~p_in[0]), .g0(~g_in[0]), .gp(node_level4_pos8_outg), .pp(node_level4_pos8_outp));
	wire node_level4_pos9_outg;
	wire node_level4_pos9_outp;
	pos_operator node_level4_pos9(.p1(node_level3_pos9_outp), .g1(node_level3_pos9_outg), .p0(node_level1_pos1_outp), .g0(node_level1_pos1_outg), .gp(node_level4_pos9_outg), .pp(node_level4_pos9_outp));
	wire node_level4_pos10_outg;
	wire node_level4_pos10_outp;
	pos_operator node_level4_pos10(.p1(node_level3_pos10_outp), .g1(node_level3_pos10_outg), .p0(~node_level2_pos2_outp), .g0(~node_level2_pos2_outg), .gp(node_level4_pos10_outg), .pp(node_level4_pos10_outp));
	wire node_level4_pos11_outg;
	wire node_level4_pos11_outp;
	pos_operator node_level4_pos11(.p1(node_level3_pos11_outp), .g1(node_level3_pos11_outg), .p0(~node_level2_pos3_outp), .g0(~node_level2_pos3_outg), .gp(node_level4_pos11_outg), .pp(node_level4_pos11_outp));
	wire node_level4_pos12_outg;
	wire node_level4_pos12_outp;
	pos_operator node_level4_pos12(.p1(node_level3_pos12_outp), .g1(node_level3_pos12_outg), .p0(node_level3_pos4_outp), .g0(node_level3_pos4_outg), .gp(node_level4_pos12_outg), .pp(node_level4_pos12_outp));
	wire node_level4_pos13_outg;
	wire node_level4_pos13_outp;
	pos_operator node_level4_pos13(.p1(node_level3_pos13_outp), .g1(node_level3_pos13_outg), .p0(node_level3_pos5_outp), .g0(node_level3_pos5_outg), .gp(node_level4_pos13_outg), .pp(node_level4_pos13_outp));
	wire node_level4_pos14_outg;
	wire node_level4_pos14_outp;
	pos_operator node_level4_pos14(.p1(node_level3_pos14_outp), .g1(node_level3_pos14_outg), .p0(node_level3_pos6_outp), .g0(node_level3_pos6_outg), .gp(node_level4_pos14_outg), .pp(node_level4_pos14_outp));
	wire node_level4_pos15_outg;
	wire node_level4_pos15_outp;
	pos_operator node_level4_pos15(.p1(node_level3_pos15_outp), .g1(node_level3_pos15_outg), .p0(node_level3_pos7_outp), .g0(node_level3_pos7_outg), .gp(node_level4_pos15_outg), .pp(node_level4_pos15_outp));
	wire node_level4_pos16_outg;
	wire node_level4_pos16_outp;
	pos_operator node_level4_pos16(.p1(node_level3_pos16_outp), .g1(node_level3_pos16_outg), .p0(node_level3_pos8_outp), .g0(node_level3_pos8_outg), .gp(node_level4_pos16_outg), .pp(node_level4_pos16_outp));
	wire node_level4_pos17_outg;
	wire node_level4_pos17_outp;
	pos_operator node_level4_pos17(.p1(node_level3_pos17_outp), .g1(node_level3_pos17_outg), .p0(node_level3_pos9_outp), .g0(node_level3_pos9_outg), .gp(node_level4_pos17_outg), .pp(node_level4_pos17_outp));
	wire node_level4_pos18_outg;
	wire node_level4_pos18_outp;
	pos_operator node_level4_pos18(.p1(node_level3_pos18_outp), .g1(node_level3_pos18_outg), .p0(node_level3_pos10_outp), .g0(node_level3_pos10_outg), .gp(node_level4_pos18_outg), .pp(node_level4_pos18_outp));
	wire node_level4_pos19_outg;
	wire node_level4_pos19_outp;
	pos_operator node_level4_pos19(.p1(node_level3_pos19_outp), .g1(node_level3_pos19_outg), .p0(node_level3_pos11_outp), .g0(node_level3_pos11_outg), .gp(node_level4_pos19_outg), .pp(node_level4_pos19_outp));
	wire node_level4_pos20_outg;
	wire node_level4_pos20_outp;
	pos_operator node_level4_pos20(.p1(node_level3_pos20_outp), .g1(node_level3_pos20_outg), .p0(node_level3_pos12_outp), .g0(node_level3_pos12_outg), .gp(node_level4_pos20_outg), .pp(node_level4_pos20_outp));
	wire node_level4_pos21_outg;
	wire node_level4_pos21_outp;
	pos_operator node_level4_pos21(.p1(node_level3_pos21_outp), .g1(node_level3_pos21_outg), .p0(node_level3_pos13_outp), .g0(node_level3_pos13_outg), .gp(node_level4_pos21_outg), .pp(node_level4_pos21_outp));
	wire node_level4_pos22_outg;
	wire node_level4_pos22_outp;
	pos_operator node_level4_pos22(.p1(node_level3_pos22_outp), .g1(node_level3_pos22_outg), .p0(node_level3_pos14_outp), .g0(node_level3_pos14_outg), .gp(node_level4_pos22_outg), .pp(node_level4_pos22_outp));
	wire node_level4_pos23_outg;
	wire node_level4_pos23_outp;
	pos_operator node_level4_pos23(.p1(node_level3_pos23_outp), .g1(node_level3_pos23_outg), .p0(node_level3_pos15_outp), .g0(node_level3_pos15_outg), .gp(node_level4_pos23_outg), .pp(node_level4_pos23_outp));
	wire node_level4_pos24_outg;
	wire node_level4_pos24_outp;
	pos_operator node_level4_pos24(.p1(node_level3_pos24_outp), .g1(node_level3_pos24_outg), .p0(node_level3_pos16_outp), .g0(node_level3_pos16_outg), .gp(node_level4_pos24_outg), .pp(node_level4_pos24_outp));
	wire node_level4_pos25_outg;
	wire node_level4_pos25_outp;
	pos_operator node_level4_pos25(.p1(node_level3_pos25_outp), .g1(node_level3_pos25_outg), .p0(node_level3_pos17_outp), .g0(node_level3_pos17_outg), .gp(node_level4_pos25_outg), .pp(node_level4_pos25_outp));
	wire node_level4_pos26_outg;
	wire node_level4_pos26_outp;
	pos_operator node_level4_pos26(.p1(node_level3_pos26_outp), .g1(node_level3_pos26_outg), .p0(node_level3_pos18_outp), .g0(node_level3_pos18_outg), .gp(node_level4_pos26_outg), .pp(node_level4_pos26_outp));
	wire node_level4_pos27_outg;
	wire node_level4_pos27_outp;
	pos_operator node_level4_pos27(.p1(node_level3_pos27_outp), .g1(node_level3_pos27_outg), .p0(node_level3_pos19_outp), .g0(node_level3_pos19_outg), .gp(node_level4_pos27_outg), .pp(node_level4_pos27_outp));
	wire node_level4_pos28_outg;
	wire node_level4_pos28_outp;
	pos_operator node_level4_pos28(.p1(node_level3_pos28_outp), .g1(node_level3_pos28_outg), .p0(node_level3_pos20_outp), .g0(node_level3_pos20_outg), .gp(node_level4_pos28_outg), .pp(node_level4_pos28_outp));
	wire node_level4_pos29_outg;
	wire node_level4_pos29_outp;
	pos_operator node_level4_pos29(.p1(node_level3_pos29_outp), .g1(node_level3_pos29_outg), .p0(node_level3_pos21_outp), .g0(node_level3_pos21_outg), .gp(node_level4_pos29_outg), .pp(node_level4_pos29_outp));
	wire node_level4_pos30_outg;
	wire node_level4_pos30_outp;
	pos_operator node_level4_pos30(.p1(node_level3_pos30_outp), .g1(node_level3_pos30_outg), .p0(node_level3_pos22_outp), .g0(node_level3_pos22_outg), .gp(node_level4_pos30_outg), .pp(node_level4_pos30_outp));
	wire node_level4_pos31_outg;
	wire node_level4_pos31_outp;
	pos_operator node_level4_pos31(.p1(node_level3_pos31_outp), .g1(node_level3_pos31_outg), .p0(node_level3_pos23_outp), .g0(node_level3_pos23_outg), .gp(node_level4_pos31_outg), .pp(node_level4_pos31_outp));
	wire node_level5_pos16_outg;
	wire node_level5_pos16_outp;
	neg_operator node_level5_pos16(.p1(node_level4_pos16_outp), .g1(node_level4_pos16_outg), .p0(p_in[0]), .g0(g_in[0]), .gp(node_level5_pos16_outg), .pp(node_level5_pos16_outp));
	wire node_level5_pos17_outg;
	wire node_level5_pos17_outp;
	neg_operator node_level5_pos17(.p1(node_level4_pos17_outp), .g1(node_level4_pos17_outg), .p0(~node_level1_pos1_outp), .g0(~node_level1_pos1_outg), .gp(node_level5_pos17_outg), .pp(node_level5_pos17_outp));
	wire node_level5_pos18_outg;
	wire node_level5_pos18_outp;
	neg_operator node_level5_pos18(.p1(node_level4_pos18_outp), .g1(node_level4_pos18_outg), .p0(node_level2_pos2_outp), .g0(node_level2_pos2_outg), .gp(node_level5_pos18_outg), .pp(node_level5_pos18_outp));
	wire node_level5_pos19_outg;
	wire node_level5_pos19_outp;
	neg_operator node_level5_pos19(.p1(node_level4_pos19_outp), .g1(node_level4_pos19_outg), .p0(node_level2_pos3_outp), .g0(node_level2_pos3_outg), .gp(node_level5_pos19_outg), .pp(node_level5_pos19_outp));
	wire node_level5_pos20_outg;
	wire node_level5_pos20_outp;
	neg_operator node_level5_pos20(.p1(node_level4_pos20_outp), .g1(node_level4_pos20_outg), .p0(~node_level3_pos4_outp), .g0(~node_level3_pos4_outg), .gp(node_level5_pos20_outg), .pp(node_level5_pos20_outp));
	wire node_level5_pos21_outg;
	wire node_level5_pos21_outp;
	neg_operator node_level5_pos21(.p1(node_level4_pos21_outp), .g1(node_level4_pos21_outg), .p0(~node_level3_pos5_outp), .g0(~node_level3_pos5_outg), .gp(node_level5_pos21_outg), .pp(node_level5_pos21_outp));
	wire node_level5_pos22_outg;
	wire node_level5_pos22_outp;
	neg_operator node_level5_pos22(.p1(node_level4_pos22_outp), .g1(node_level4_pos22_outg), .p0(~node_level3_pos6_outp), .g0(~node_level3_pos6_outg), .gp(node_level5_pos22_outg), .pp(node_level5_pos22_outp));
	wire node_level5_pos23_outg;
	wire node_level5_pos23_outp;
	neg_operator node_level5_pos23(.p1(node_level4_pos23_outp), .g1(node_level4_pos23_outg), .p0(~node_level3_pos7_outp), .g0(~node_level3_pos7_outg), .gp(node_level5_pos23_outg), .pp(node_level5_pos23_outp));
	wire node_level5_pos24_outg;
	wire node_level5_pos24_outp;
	neg_operator node_level5_pos24(.p1(node_level4_pos24_outp), .g1(node_level4_pos24_outg), .p0(node_level4_pos8_outp), .g0(node_level4_pos8_outg), .gp(node_level5_pos24_outg), .pp(node_level5_pos24_outp));
	wire node_level5_pos25_outg;
	wire node_level5_pos25_outp;
	neg_operator node_level5_pos25(.p1(node_level4_pos25_outp), .g1(node_level4_pos25_outg), .p0(node_level4_pos9_outp), .g0(node_level4_pos9_outg), .gp(node_level5_pos25_outg), .pp(node_level5_pos25_outp));
	wire node_level5_pos26_outg;
	wire node_level5_pos26_outp;
	neg_operator node_level5_pos26(.p1(node_level4_pos26_outp), .g1(node_level4_pos26_outg), .p0(node_level4_pos10_outp), .g0(node_level4_pos10_outg), .gp(node_level5_pos26_outg), .pp(node_level5_pos26_outp));
	wire node_level5_pos27_outg;
	wire node_level5_pos27_outp;
	neg_operator node_level5_pos27(.p1(node_level4_pos27_outp), .g1(node_level4_pos27_outg), .p0(node_level4_pos11_outp), .g0(node_level4_pos11_outg), .gp(node_level5_pos27_outg), .pp(node_level5_pos27_outp));
	wire node_level5_pos28_outg;
	wire node_level5_pos28_outp;
	neg_operator node_level5_pos28(.p1(node_level4_pos28_outp), .g1(node_level4_pos28_outg), .p0(node_level4_pos12_outp), .g0(node_level4_pos12_outg), .gp(node_level5_pos28_outg), .pp(node_level5_pos28_outp));
	wire node_level5_pos29_outg;
	wire node_level5_pos29_outp;
	neg_operator node_level5_pos29(.p1(node_level4_pos29_outp), .g1(node_level4_pos29_outg), .p0(node_level4_pos13_outp), .g0(node_level4_pos13_outg), .gp(node_level5_pos29_outg), .pp(node_level5_pos29_outp));
	wire node_level5_pos30_outg;
	wire node_level5_pos30_outp;
	neg_operator node_level5_pos30(.p1(node_level4_pos30_outp), .g1(node_level4_pos30_outg), .p0(node_level4_pos14_outp), .g0(node_level4_pos14_outg), .gp(node_level5_pos30_outg), .pp(node_level5_pos30_outp));
	wire node_level5_pos31_outg;
	wire node_level5_pos31_outp;
	neg_operator node_level5_pos31(.p1(node_level4_pos31_outp), .g1(node_level4_pos31_outg), .p0(node_level4_pos15_outp), .g0(node_level4_pos15_outg), .gp(node_level5_pos31_outg), .pp(node_level5_pos31_outp));


	assign s[0] = p_in[0] ^ cin;
	assign s[1] = p_in[1] ^ g_in[0];
	assign s[2] = p_in[2] ^ ~node_level1_pos1_outg;
	assign s[3] = p_in[3] ^ node_level2_pos2_outg;
	assign s[4] = p_in[4] ^ node_level2_pos3_outg;
	assign s[5] = p_in[5] ^ ~node_level3_pos4_outg;
	assign s[6] = p_in[6] ^ ~node_level3_pos5_outg;
	assign s[7] = p_in[7] ^ ~node_level3_pos6_outg;
	assign s[8] = p_in[8] ^ ~node_level3_pos7_outg;
	assign s[9] = p_in[9] ^ node_level4_pos8_outg;
	assign s[10] = p_in[10] ^ node_level4_pos9_outg;
	assign s[11] = p_in[11] ^ node_level4_pos10_outg;
	assign s[12] = p_in[12] ^ node_level4_pos11_outg;
	assign s[13] = p_in[13] ^ node_level4_pos12_outg;
	assign s[14] = p_in[14] ^ node_level4_pos13_outg;
	assign s[15] = p_in[15] ^ node_level4_pos14_outg;
	assign s[16] = p_in[16] ^ node_level4_pos15_outg;
	assign s[17] = p_in[17] ^ ~node_level5_pos16_outg;
	assign s[18] = p_in[18] ^ ~node_level5_pos17_outg;
	assign s[19] = p_in[19] ^ ~node_level5_pos18_outg;
	assign s[20] = p_in[20] ^ ~node_level5_pos19_outg;
	assign s[21] = p_in[21] ^ ~node_level5_pos20_outg;
	assign s[22] = p_in[22] ^ ~node_level5_pos21_outg;
	assign s[23] = p_in[23] ^ ~node_level5_pos22_outg;
	assign s[24] = p_in[24] ^ ~node_level5_pos23_outg;
	assign s[25] = p_in[25] ^ ~node_level5_pos24_outg;
	assign s[26] = p_in[26] ^ ~node_level5_pos25_outg;
	assign s[27] = p_in[27] ^ ~node_level5_pos26_outg;
	assign s[28] = p_in[28] ^ ~node_level5_pos27_outg;
	assign s[29] = p_in[29] ^ ~node_level5_pos28_outg;
	assign s[30] = p_in[30] ^ ~node_level5_pos29_outg;
	assign s[31] = p_in[31] ^ ~node_level5_pos30_outg;
	assign cout = (x1[31] & x2[31]) | (~s[31] & (x1[31] | x2[31]));
endmodule
